`timescale 1ns / 1ps

// ---------------------------------------------------------------------
// UDP����ģ�� 
// ---------------------------------------------------------------------


module udp_tx(
    input                   clk,
    input                   rst,

    input                   tx_start_en,                // ����UDP����ʹ���ź�
    input           [15:0]  tx_byte_num,                // ����UDP�������ݶ��ֽ���
    input           [7:0]   tx_data,                    // UDP���ݶ������ֽ�
    input           [31:0]  crc_data,
    input           [7:0]   crc_next,
    input           [31:0]  des_ip,
    input           [47:0]  des_mac,

    output  reg             crc_clr,
    output  reg             crc_en,
    output  reg             gmii_tx_en,                 // ����gmii����ʹ���ź�
    output  reg     [7:0]   gmii_txd,
    output  reg             tx_done,                    // ����UDP���ݱ�������ź�s
    output  reg             tx_req 
    );

    // parameter define
    parameter   BOARD_MAC  = 48'h00_11_22_33_44_55;
    parameter   BOARD_IP   = {8'd192, 8'd168, 8'd0, 8'd2};
    parameter   DES_MAC    = 48'hff_ff_ff_ff_ff_ff;
    parameter   DES_IP     = {8'd192,8'd168,8'd0,8'd3}; 

    localparam  ETH_TYPE        = 16'h0800;                 // �ϲ�Э��ΪIP����
    localparam  MIN_DATA_NUM    = 16'd18;                   // UDP�������ݲ�����С���ȣ�46-20(IPͷ������)-8(UDPͷ������)
    localparam  UDP_TYPE        = 8'd17;                    // UDPЭ���17

    localparam  st_idle         = 7'b000_0001;
    localparam  st_check_ip     = 7'b000_0010;              // ����IPͷ��У���
    localparam  st_preamble     = 7'b000_0100;
    localparam  st_eth_header   = 7'b000_1000;
    localparam  st_ip_header    = 7'b001_0000;              // ����20�ֽ�IPͷ��8�ֽ�UDPͷ
    localparam  st_tx_data      = 7'b010_0000;
    localparam  st_crc          = 7'b100_0000;

    // reg define
    reg [6:0]   cur_state;
    reg [6:0]   next_state;
    reg [7:0]   preamble[7:0];
    reg [7:0]   eth_header[13:0];
    reg [31:0]  ip_header[6:0];                             // IPͷ+UDPͷ��28��
    reg         start_en_d0;
    reg         start_en_d1;
    reg         start_en_d2;                                // ��tx_start_en�źŴ�����
    reg         trig_tx_en;                                 // ������ʼ�����ź�
    reg [15:0]  tx_data_num;                                // �Ĵ����ݶ��ֽ���
    reg [15:0]  total_num;                                  // IP���ĵ����ֽ���
    reg [15:0]  udp_num;                                    // UDP���ĵ����ֽ���
    reg         skip_en;
    reg [4:0]   cnt;
    reg [31:0]  check_buffer;                               // IPͷУ��ͼ��㻺��
    reg [1:0]   tx_byte_sel;                                 // 4�ֽڷ��ͼ�����
    reg [15:0]  data_cnt;                                   // ���ݶ��ֽڼ���ָ��
    reg         tx_done_t;
    reg [15:0]  real_add_cnt;                               // ʵ����Ҫ�����ֽ��������ĳ���С��48�ֽ�ʱ��

    // wire define
    wire            pos_start_en;                           // tx_start_en��������
    wire    [15:0]  real_tx_data_num;                       // ʵ�ʷ��͵��ֽ�����������̫�������ֽ�Ҫ��

    assign  pos_start_en = ~start_en_d2 & start_en_d1;
    assign  real_tx_data_num = (tx_data_num >= MIN_DATA_NUM) ? tx_data_num : MIN_DATA_NUM;

    // �����Ĳɼ�tx_start_en��������
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            start_en_d0 <= 1'b0;
            start_en_d1 <= 1'b0;
            start_en_d2 <= 1'b0;
        end
        else begin
            start_en_d0 <= tx_start_en;
            start_en_d1 <= start_en_d0;
            start_en_d2 <= start_en_d1;
        end
    end

    // �Ĵ�UDP���ݶγ���
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            tx_data_num <= 16'd0;
            total_num   <= 16'd0;
            udp_num     <= 16'd0;
        end
        else begin
            if(pos_start_en && (cur_state == st_idle)) begin
                tx_data_num <= tx_byte_num;                     // �Ĵ�UDP�����ֶγ���
                udp_num     <= tx_byte_num + 16'd8;
                total_num   <= tx_byte_num + 16'd28;            // �ܳ��ȣ�UDP���ݶγ���+IPͷ(20)+UDPͷ����(8)
            end
        end
    end

    // �Ĵ�һ�Ĵ��������źţ�Ϊ����������ݶγ��Ⱥ��ܳ��ȵļĴ�
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            trig_tx_en <= 1'b0;
        end
        else begin
            trig_tx_en <= pos_start_en;
        end
    end

    // ---------------------------  ����UDP����״̬��   ----------------------------
    always @(posedge clk or posedge rst) begin
        if(rst)
            cur_state <= st_idle;
        else
            cur_state <= next_state;
    end

    always @(*) begin
        next_state = st_idle;
        case(cur_state)
            st_idle:begin
                if(skip_en)
                    next_state = st_check_ip;
                else
                    next_state = st_idle;
            end

            st_check_ip:begin
                if(skip_en)
                    next_state = st_preamble;
                else
                    next_state = st_check_ip;
            end

            st_preamble:begin
                if(skip_en)
                    next_state = st_eth_header;
                else
                    next_state = st_preamble;
            end

            st_eth_header:begin
                if(skip_en)
                    next_state = st_ip_header;
                else
                    next_state = st_eth_header;
            end

            st_ip_header:begin
                if(skip_en)
                    next_state = st_tx_data;
                else
                    next_state =st_ip_header;
            end

            st_tx_data:begin
                if(skip_en)
                    next_state = st_crc;
                else    
                    next_state = st_tx_data;
            end

            st_crc:begin
                if(skip_en)
                    next_state = st_idle;
                else
                    next_state = st_crc;
            end

            default:next_state = st_idle;
        endcase
    end

    always @(posedge clk or posedge rst) begin
        if(rst) begin
            // �Ĵ�����ʼ��
            skip_en                 <= 1'b0; 
            cnt                     <= 5'd0;
            check_buffer            <= 32'd0;
            ip_header[1][31:16]     <= 16'd0;
            tx_byte_sel             <= 2'd0;
            crc_en                  <= 1'b0;
            gmii_tx_en              <= 1'b0;
            gmii_txd                <= 8'd0;
            tx_req                  <= 1'b0;
            tx_done_t               <= 1'b0; 
            data_cnt                <= 16'd0;
            real_add_cnt            <= 5'd0;

            //ǰ���� 7��8'h55 + 1��8'hd5 
            preamble[0] <= 8'h55;                
            preamble[1] <= 8'h55;
            preamble[2] <= 8'h55;
            preamble[3] <= 8'h55;
            preamble[4] <= 8'h55;
            preamble[5] <= 8'h55;
            preamble[6] <= 8'h55;
            preamble[7] <= 8'hd5;

            // ��̫ͷ
            eth_header[0] <= DES_MAC[47:40];            // Ŀ��mac
            eth_header[1] <= DES_MAC[39:32];
            eth_header[2] <= DES_MAC[31:24];
            eth_header[3] <= DES_MAC[23:16];
            eth_header[4] <= DES_MAC[15:8];
            eth_header[5] <= DES_MAC[7:0];

            eth_header[6] <= BOARD_MAC[47:40];          // ���ͷ�mac
            eth_header[7] <= BOARD_MAC[39:32];
            eth_header[8] <= BOARD_MAC[31:24];
            eth_header[9] <= BOARD_MAC[23:16];
            eth_header[10] <= BOARD_MAC[15:8];
            eth_header[11] <= BOARD_MAC[7:0];

            eth_header[12] <= ETH_TYPE[15:8];           // ��̫����
            eth_header[13] <= ETH_TYPE[7:0];

        end
        else begin
            skip_en <= 1'b0;
            tx_done_t <= 1'b0;
            gmii_tx_en <= 1'b0;
            crc_en <= 1'b0;
            case(next_state)
                st_idle:begin
                    if(trig_tx_en) begin
                        skip_en <= 1'b1;
                        // �汾�ţ�4���ײ����ȣ�5����λ��4bytes����20�ֽڣ�,��������00���ܳ���
                        ip_header[0] <= {8'h45, 8'h00, total_num};
                        // 16λ���ı�ʶ����ͬһ�������з�Ƭ��ʶ����ͬ
                        ip_header[1][31:16] <= ip_header[1][31:16] + 16'd1;             // ÿ����һ�Σ���ʶ����1
                        // ��־��Ƭƫ�ƣ�010����Ƭ��Ƭƫ��Ϊ0
                        ip_header[1][15:0]  <= 16'h4000;                                // ��ʹ�÷�Ƭ
                        // ����ʱ�䣬Э�����ͣ�80����ʱ��128��Э������17��UDP���ײ�У�����ʹ��0
                        ip_header[2] <= {8'h80, UDP_TYPE, 16'h0000};
                        // ԴIP��ַ
                        ip_header[3] <= BOARD_IP;
                        // Ŀ��IP��ַ
                        if(des_ip != 32'd0)
                            ip_header[4] <= des_ip;
                        else
                            ip_header[4] <= DES_IP;
                        // UDPͷ
                        // Դ�˿���Ŀ�Ķ˿�
                        ip_header[5] <= {16'd1234, 16'd1234};                           // Դ�˿ں�Ŀ�Ķ˿ھ�Ϊ1234
                        // UDP���Ⱥ�У��ͣ���ʹ�ã�Ĭ��Ϊ0��
                        ip_header[6] <= {udp_num, 16'd0};
                        
                        // ������̫ͷ�е�Ŀ��mac
                        if(des_mac != 48'd0) begin
                            eth_header[0]  <= des_mac[47:40];
                            eth_header[1]  <= des_mac[39:32];
                            eth_header[2]  <= des_mac[31:24];
                            eth_header[3]  <= des_mac[23:16];
                            eth_header[4]  <= des_mac[15:8] ;
                            eth_header[5]  <= des_mac[7:0]  ;
                        end
                    end
                end

                st_check_ip:begin
                    cnt <= cnt + 5'd1;
                    if(cnt == 5'd0) begin
                        check_buffer <= ip_header[0][31:16] + ip_header[0][15:0]
                                        + ip_header[1][31:16] + ip_header[1][15:0]
                                        + ip_header[2][31:16] + ip_header[2][15:0]
                                        + ip_header[3][31:16] + ip_header[3][15:0]
                                        + ip_header[4][31:16] + ip_header[4][15:0];
                    end
                    else if(cnt == 5'd1) begin
                        check_buffer <= check_buffer[31:16] + check_buffer[15:0];       // check_buffer��32λ��
                    end
                    else if(cnt == 5'd2) begin
                        check_buffer <= check_buffer[31:16] + check_buffer[15:0];       //�����ٴγ��ֽ�λ����һ��
                    end             
                    else if(cnt == 5'd3) begin
                        skip_en <= 1'b1;
                        cnt <= 5'd0;
                        ip_header[2][15:0] <= ~check_buffer[15:0];
                    end
                end

                st_preamble:begin
                    gmii_tx_en <= 1'b1;
                    gmii_txd <= preamble[cnt];
                    if(cnt == 5'd7) begin
                        skip_en <= 1'b1;
                        cnt <= 5'd0;
                    end
                    else 
                        cnt <= cnt + 5'd1;
                end

                st_eth_header:begin
                    gmii_tx_en <= 1'b1;
                    crc_en <= 1'b1;
                    gmii_txd <= eth_header[cnt];
                    if(cnt == 5'd13) begin
                        skip_en <= 1'b1;
                        cnt <= 5'd0;
                    end
                    else
                        cnt <= cnt + 5'd1;
                end

                st_ip_header:begin
                    gmii_tx_en <= 1'b1;
                    crc_en <= 1'b1;
                    tx_byte_sel <= tx_byte_sel + 2'd1;
                    // ˫��ѭ������
                    if(tx_byte_sel == 2'd0)
                        gmii_txd <= ip_header[cnt][31:24];
                    else if(tx_byte_sel == 2'd1)
                        gmii_txd <= ip_header[cnt][23:16];
                    else if(tx_byte_sel == 2'd2) begin
                        gmii_txd <= ip_header[cnt][15:8];
                        if(cnt == 5'd6) 
                            // ��ǰ�������ݣ��ȴ���Ч�źŵ���ʱֱ�ӷ���
                            tx_req <= 1'b1;
                    end
                    else if(tx_byte_sel == 2'd3) begin
                        gmii_txd <= ip_header[cnt][7:0];
                        if(cnt == 5'd6) begin
                            skip_en <= 1'b1;
                            cnt <= 5'd0;
                            
                        end
                        else
                            cnt <= cnt + 5'd1;
                    end
                end

                st_tx_data:begin
                    gmii_tx_en <= 1'b1;
                    crc_en <= 1'b1;
                    tx_byte_sel <= 2'd0;
                    gmii_txd <= tx_data;

                    if(data_cnt < tx_data_num - 16'd1)
                        data_cnt <= data_cnt + 16'd1;
                    else if(data_cnt == tx_data_num - 16'd1) begin
                        if(data_cnt + real_add_cnt < real_tx_data_num - 16'd1)
                            real_add_cnt <= real_add_cnt + 16'd1;       // ������Ҫ�������ֽ�
                        else begin
                            skip_en <= 1'b1;
                            data_cnt <= 16'd0;
                            real_add_cnt <= 16'd0;
                        end
                    end

                    if(data_cnt == tx_data_num - 16'd2) 
                        tx_req <= 1'b0;

                end

                st_crc:begin
                    gmii_tx_en <= 1'b1;
                    tx_byte_sel <= tx_byte_sel + 2'd1;

                    if(tx_byte_sel == 2'd0)
                        gmii_txd <= {~crc_next[0], ~crc_next[1], ~crc_next[2],~crc_next[3],
                                    ~crc_next[4], ~crc_next[5], ~crc_next[6],~crc_next[7]};
                    else if(tx_byte_sel == 2'd1)
                        gmii_txd <= {~crc_data[16], ~crc_data[17], ~crc_data[18],~crc_data[19],
                                    ~crc_data[20], ~crc_data[21], ~crc_data[22],~crc_data[23]};
                    else if(tx_byte_sel == 2'd2) begin
                        gmii_txd <= {~crc_data[8], ~crc_data[9], ~crc_data[10],~crc_data[11],
                                    ~crc_data[12], ~crc_data[13], ~crc_data[14],~crc_data[15]};                              
                    end
                    else if(tx_byte_sel == 2'd3) begin
                        gmii_txd <= {~crc_data[0], ~crc_data[1], ~crc_data[2],~crc_data[3],
                                    ~crc_data[4], ~crc_data[5], ~crc_data[6],~crc_data[7]};  
                        tx_done_t <= 1'b1;
                        skip_en <= 1'b1;
                    end     
                end

                default: ;
            endcase
        end
    end

    //��������źż�crcֵ��λ�ź�
    always @(posedge clk or negedge rst) begin
        if(rst) begin
            tx_done <= 1'b0;
            crc_clr <= 1'b0;
        end
        else begin
            tx_done <= tx_done_t;
            crc_clr <= tx_done_t;
        end
    end


endmodule
