`timescale 1ns / 1ps

module tb_arp_top();

// ====================== ʱ�Ӻ͸�λ�ź� ======================
reg sys_clk_p;
reg sys_clk_n;

reg gtrefclk_p;
reg gtrefclk_n;

reg sys_rst_n;

// ʱ�Ӳ���
parameter SYS_CLK_PERIOD = 5;     // 200MHz (5ns����)
parameter GTREFCLK_PERIOD = 8;    // 125MHz (8ns����)

// ʱ������
initial begin
    sys_clk_p = 1'b0;
    forever #(SYS_CLK_PERIOD/2) sys_clk_p = ~sys_clk_p;
end

assign sys_clk_n = ~sys_clk_p;

initial begin
    gtrefclk_p = 1'b0;
    forever #(GTREFCLK_PERIOD/2) gtrefclk_p = ~gtrefclk_p;
end

assign gtrefclk_n = ~gtrefclk_p;

// ====================== ��λ���� ======================
initial begin
    sys_rst_n = 1'b0;
    #100 sys_rst_n = 1'b1;  // 100ns���ͷŸ�λ
end

// ====================== ʵ����DUT ======================
wire txp, txn;
wire phy_rst_n;
wire led_link;

// ����ARP��������
wire [7:0] gmii_tx_data;
wire gmii_tx_en;
wire gmii_tx_err;

// �޸�test_top������ڲ�GMII�ź�������֤
test_top dut (
    .sys_clk_p(sys_clk_p),
    .sys_clk_n(sys_clk_n),
    .gtrefclk_p(gtrefclk_p),
    .gtrefclk_n(gtrefclk_n),
    .sys_rst_n(sys_rst_n),
    .phy_rst_n(phy_rst_n),
    
    // SGMII�ӿ� - ���ӵ�����PHY
    .txp(txp),
    .txn(txn),
    .rxp(1'b0),  // ���ղ����գ���Ϊ����ֻ���Է���
    .rxn(1'b1),
    
    // ״ָ̬ʾ
    .led_link(led_link),
    
    // ���ڲ��Ե��ڲ��źţ���Ҫ��test_top������Ϊ�����
    .test_gmii_tx_data(gmii_tx_data),
    .test_gmii_tx_en(gmii_tx_en),
    .test_gmii_tx_err(gmii_tx_err)
);

// ====================== ����PHY������ ======================
// ���ڲ������֤ARP���ݰ�
reg [7:0] packet_buffer [0:511];
reg [9:0] packet_index = 0;
reg packet_capturing = 0;
reg [31:0] byte_counter = 0;

// ����GMII������
always @(posedge gmii_clk) begin
    if (!sys_rst_n) begin
        packet_index <= 0;
        packet_capturing <= 0;
        byte_counter <= 0;
    end else begin
        byte_counter <= byte_counter + 1;
        
        // ���֡��ʼ��ǰ����+SFD��
        if (gmii_tx_en && gmii_tx_data == 8'hD5 && packet_index == 7) begin
            packet_capturing <= 1;
            packet_index <= 0;
            $display("[%0t] INFO: Start of Frame Detected", $time);
        end 
        // ����֡����
        else if (gmii_tx_en && packet_capturing) begin
            packet_buffer[packet_index] <= gmii_tx_data;
            packet_index <= packet_index + 1;
            
            // ��֡������⣨��ʵ����Ӧ�ü��IFG��
            if (packet_index > 100) begin
                packet_capturing <= 0;
                $display("[%0t] INFO: Frame captured, length = %0d bytes", $time, packet_index);
                verify_arp_packet();
            end
        end
        // ֡����
        else if (!gmii_tx_en && packet_capturing) begin
            packet_capturing <= 0;
            $display("[%0t] INFO: End of Frame, captured %0d bytes", $time, packet_index);
            verify_arp_packet();
        end
    end
end

// ====================== ARP���ݰ���֤ ======================
task verify_arp_packet;
    integer i;
    reg [47:0] dest_mac;
    reg [47:0] src_mac;
    reg [15:0] eth_type;
    reg [15:0] arp_hw_type;
    reg [15:0] arp_protocol;
    reg [7:0] arp_hw_len;
    reg [7:0] arp_prot_len;
    reg [15:0] arp_opcode;
    reg [47:0] arp_src_mac;
    reg [31:0] arp_src_ip;
    reg [47:0] arp_dest_mac;
    reg [31:0] arp_dest_ip;
begin
    $display("\n========== ARP Packet Verification ==========");
    
    // ��֤��̫��ͷ������SFD֮��ʼ��
    dest_mac = {packet_buffer[0], packet_buffer[1], packet_buffer[2], 
                packet_buffer[3], packet_buffer[4], packet_buffer[5]};
    src_mac = {packet_buffer[6], packet_buffer[7], packet_buffer[8], 
               packet_buffer[9], packet_buffer[10], packet_buffer[11]};
    eth_type = {packet_buffer[12], packet_buffer[13]};
         
    $display("Destination MAC: %02x:%02x:%02x:%02x:%02x:%02x",
             dest_mac[47:40], dest_mac[39:32], dest_mac[31:24],
             dest_mac[23:16], dest_mac[15:8], dest_mac[7:0]);
    $display("Source MAC: %02x:%02x:%02x:%02x:%02x:%02x",
             src_mac[47:40], src_mac[39:32], src_mac[31:24],
             src_mac[23:16], src_mac[15:8], src_mac[7:0]);
    $display("EtherType: 0x%04x", eth_type);
    
    // ��֤ARP���ݲ���
    arp_hw_type = {packet_buffer[14], packet_buffer[15]};
    arp_protocol = {packet_buffer[16], packet_buffer[17]};
    arp_hw_len = packet_buffer[18];
    arp_prot_len = packet_buffer[19];
    arp_opcode = {packet_buffer[20], packet_buffer[21]};
    arp_src_mac = {packet_buffer[22], packet_buffer[23], packet_buffer[24],
                   packet_buffer[25], packet_buffer[26], packet_buffer[27]};
    arp_src_ip = {packet_buffer[28], packet_buffer[29], 
                  packet_buffer[30], packet_buffer[31]};
    arp_dest_mac = {packet_buffer[32], packet_buffer[33], packet_buffer[34],
                    packet_buffer[35], packet_buffer[36], packet_buffer[37]};
    arp_dest_ip = {packet_buffer[38], packet_buffer[39],
                   packet_buffer[40], packet_buffer[41]};
    
    $display("\nARP Header:");
    $display("  HW Type: 0x%04x (1=Ethernet)", arp_hw_type);
    $display("  Protocol: 0x%04x (0x0800=IPv4)", arp_protocol);
    $display("  HW Addr Len: %0d", arp_hw_len);
    $display("  Protocol Addr Len: %0d", arp_prot_len);
    $display("  Opcode: 0x%04x (1=Request, 2=Reply)", arp_opcode);
    $display("  Sender MAC: %02x:%02x:%02x:%02x:%02x:%02x",
             arp_src_mac[47:40], arp_src_mac[39:32], arp_src_mac[31:24],
             arp_src_mac[23:16], arp_src_mac[15:8], arp_src_mac[7:0]);
    $display("  Sender IP: %0d.%0d.%0d.%0d",
             arp_src_ip[31:24], arp_src_ip[23:16], arp_src_ip[15:8], arp_src_ip[7:0]);
    $display("  Target MAC: %02x:%02x:%02x:%02x:%02x:%02x",
             arp_dest_mac[47:40], arp_dest_mac[39:32], arp_dest_mac[31:24],
             arp_dest_mac[23:16], arp_dest_mac[15:8], arp_dest_mac[7:0]);
    $display("  Target IP: %0d.%0d.%0d.%0d",
             arp_dest_ip[31:24], arp_dest_ip[23:16], arp_dest_ip[15:8], arp_dest_ip[7:0]);
    
    // ��֤����ֵ
    if (dest_mac == 48'hFFFFFFFFFFFF) begin
        $display("\n? Destination MAC is broadcast (correct)");
    end else begin
        $display("\n? Destination MAC error: expected broadcast");
    end
    
    if (src_mac == 48'h000A3501FEC0) begin
        $display("? Source MAC matches expected value");
    end else begin
        $display("? Source MAC error: expected 00:0A:35:01:FE:C0");
    end
    
    if (eth_type == 16'h0806) begin
        $display("? EtherType is ARP (0x0806)");
    end else begin
        $display("? EtherType error: expected 0x0806");
    end
    
    if (arp_opcode == 16'h0001) begin
        $display("? ARP Opcode is Request (0x0001)");
    end else begin
        $display("? ARP Opcode error: expected 0x0001");
    end
    
    if (arp_dest_ip == 32'hC0A80003) begin
        $display("? Target IP is 192.168.0.3");
    end else begin
        $display("? Target IP error: expected 192.168.0.3");
    end
    
    // ��֤CRC�����4�ֽڣ�
    $display("\nFrame CRC (last 4 bytes):");
    for (i = packet_index-4; i < packet_index; i = i+1) begin
        $write("0x%02x ", packet_buffer[i]);
    end
    $display("");
    
    $display("============================================\n");
end
endtask

// ====================== GMIIʱ�� ======================
wire gmii_clk;
// ��DUT�л�ȡuserclk2��GMIIʱ�ӣ�
assign gmii_clk = dut.userclk2;

// ====================== �źż�� ======================
// ��عؼ�״̬�ź�
initial begin
    $timeformat(-9, 3, " ns", 10);
    $display("\n========== ARP���Ͳ��Կ�ʼ ==========");
    
    // �ȴ�ϵͳ�ȶ�
    wait(sys_rst_n == 1'b1);
    $display("[%0t] INFO: System reset released", $time);
    
    // �ȴ�PCS/PMA��λ���
    wait(dut.resetdone == 1'b1);
    $display("[%0t] INFO: PCS/PMA reset done", $time);
    
    // �ȴ�ARPģ�鸴λ���
    #2000000; // �ȴ�2msȷ��ARPģ�鸴λ���
    
    $display("[%0t] INFO: Waiting for ARP packet transmission...", $time);
    
    // ���GMII�����ź�
    fork
        // ���֡��ʼ
        begin
            @(posedge gmii_tx_en);
            $display("[%0t] INFO: GMII TX_EN asserted, ARP transmission started", $time);
        end
        
        // ��ʱ���
        begin
            #20000000; // �ȴ�20ms
            if (packet_index == 0) begin
                $display("[%0t] ERROR: No ARP packet detected within timeout!", $time);
                $finish;
            end
        end
        
        // ��ض��ARP��
        begin
            repeat(3) begin  // ���3��ARP��
                wait(packet_index > 50);
                #1000;
                packet_index = 0;  // ���ü�����׼����һ����
                $display("[%0t] INFO: Waiting for next ARP packet...", $time);
            end
            $display("\n[%0t] INFO: Successfully verified 3 ARP packets", $time);
            #10000;
            $finish;
        end
    join
    
end

// ====================== ������� ======================
initial begin
    // ����VCD�ļ����ڲ��β鿴
    $dumpfile("arp_test.vcd");
    $dumpvars(0, tb_arp_top);
    
    // ����ʹ��FSDB�����֧�֣�
    // $fsdbDumpfile("arp_test.fsdb");
    // $fsdbDumpvars(0, tb_arp_top);
end

// ====================== ���Լ��� ======================
// ��������Ӷ���Ĳ��Լ��������磺
// 1. ģ��PHY״̬�仯
// 2. ���Բ�ͬ��ARP����
// 3. ���Դ���ע��

// ģ���źż��
reg signal_detect = 1'b1;
initial begin
    #5000000 signal_detect = 1'b0;  // 5us��ģ���źŶ�ʧ
    #200000 signal_detect = 1'b1;   // 200ns��ָ��ź�
end

endmodule