`timescale 1ns / 1ps

// --------------------------------------------------------
// icmp���ݱ��Ľ����߼�
// ���ڻظ�����pingӦ������
// --------------------------------------------------------

module icmp_rx(
    input                       gmii_rx_clk,
    input                       gmii_rx_dv,
    input               [7:0]   gmii_rxd,
    input                       rst,

    output   reg        [15:0]  icmp_id,                    // icmp��id�ţ���ͬid��ʾһ��icmpӦ��
    output   reg        [15:0]  icmp_seq,                   // icmp���кţ���ʶicmp���ĵ�����
    output   reg        [15:0]  rec_byte_num,               // ����icmp����payload���ֽ���
    output   reg        [7:0]   rec_data,                   // icmp���ĵ����ݣ����뵽FIFO��
    output   reg        [31:0]  reply_check_sum,            // ͷ��У���
    output   reg                rec_en,                     // ����icmp����ʹ�ܣ�����FIFO������ʹ��
    output   reg                rec_pkt_done                // �������ݰ����
    );

    // parameter define
    parameter BOARD_MAC = 48'h00_11_22_33_44_55;
    parameter BOARD_IP  = {8'd192, 8'd168, 8'd0, 8'd2};

    // ״̬������
    localparam st_idle              = 7'b000_0001;
    localparam st_preamble          = 7'b000_0010;
    localparam st_eth_header        = 7'b000_0100;
    localparam st_ip_header         = 7'b000_1000;
    localparam st_icmp_header       = 7'b001_0000;
    localparam st_rx_data           = 7'b010_0000;
    localparam st_rx_end            = 7'b100_0000;

    // ��̫�����Ͷ���
    localparam ETH_TYPE     = 16'h0800;         // ��̫��Э�����ͣ�IP
    localparam ICMP_TYPE    = 8'd1;             // ICMPЭ������

    // ICMP��������
    localparam ECHO_REQUEST = 8'h08;            // ICMP���������ǻ�������

    // reg define
    reg [6:0]   cur_state;
    reg [6:0]   next_state;
    reg         skip_en;
    reg         error_en;
    reg [4:0]   cnt;
    reg [47:0]  des_mac;                        // ICMP�Ƕ�����arp����һ�ֱ��ģ������ڸ���
    reg [31:0]  des_ip;
    reg [15:0]  eth_type;                       // ��̫������
    reg [5:0]   ip_head_byte_num;               // ipͷ�������ֽڼ���
    reg [15:0]  ip_total_length;                // IP�����ܳ���
    reg [1:0]   rec_en_cnt;                     // 8bitת32bit������
    reg [7:0]   icmp_type;                      // ICMP�������ͣ����ڱ�ʶ����Ĳ���Ļ��߲�ѯ���͵ı��汨��
    reg [7:0]   icmp_code;                      // ICMP���Ĵ��룺����ICMP����ĵ����ͣ���һ�����������ԭ��

    reg [15:0]  icmp_checksum;                   // ��������ͷ��У���
    reg [15:0]  icmp_data_length;                // ICMP��Ч�����ܳ���
    reg [15:0]  icmp_rx_cnt;                     // ICMP���������ֽڼ�����
    reg [7:0]   icmp_rx_data_d0;                 // ����һ��icmp���ݣ�ͷ��У���16bit����һ��
    reg [31:0]  reply_checksum_add;              // ͷ��У��ͼӷ���


// ------------------------------ICMP�������ݴ���״̬��----------------------------------
    always @(posedge gmii_rx_clk or posedge rst) begin
        if(rst)
            cur_state <= st_idle;
        else
            cur_state <= next_state;
    end

    always @(*) begin
        next_state = st_idle;
        case(cur_state)
            st_idle:begin
                if(skip_en)
                    next_state = st_preamble;
                else
                    next_state = st_idle;
            end

            st_preamble:begin
                if(skip_en)
                    next_state = st_eth_header;
                else if(error_en)
                    next_state = st_rx_end;
                else
                    next_state = st_preamble;
            end

            st_eth_header:begin
                if(skip_en)
                    next_state = st_ip_header;
                else if(error_en)
                    next_state = st_rx_end;
                else
                    next_state = st_eth_header;
            end

            st_ip_header:begin
                if(skip_en)
                    next_state = st_icmp_header;
                else if(error_en)
                    next_state = st_rx_end;
                else
                    next_state = st_ip_header;
            end

            st_icmp_header:begin
                if(skip_en)
                    next_state = st_rx_data;
                else if(error_en)
                    next_state = st_rx_end;
                else
                    next_state = st_icmp_header;
            end

            st_rx_data:begin
                if(skip_en)
                    next_state = st_rx_end;
                else
                    next_state = st_rx_data;
            end

            st_rx_end:begin
                if(skip_en)
                    next_state = st_idle;
                else
                    next_state = st_rx_end;
            end

            default: next_state = st_idle;
        endcase
    end

    always @(posedge gmii_rx_clk or posedge rst) begin
        if(rst) begin
            skip_en                 <= 1'd0;
            error_en                <= 1'd0;
            cnt                     <= 5'd0;
            des_mac                 <= 48'd0;
            des_ip                  <= 32'd0;
            eth_type                <= 16'd0;
            ip_head_byte_num        <= 6'd0;
            ip_total_length         <= 16'd0;
            rec_en_cnt              <= 2'd0;
            icmp_type               <= 8'd0;
            icmp_code               <= 8'd0;
            icmp_checksum           <= 16'd0;
            icmp_data_length        <= 16'd0;
            icmp_rx_cnt             <= 16'd0;
            icmp_rx_data_d0         <= 8'd0;
            reply_checksum_add      <= 32'd0;
            icmp_id                 <= 16'd0;  
            icmp_seq                <= 16'd0;
            rec_byte_num            <= 16'd0;
            rec_data                <= 8'd0;
            reply_check_sum         <= 32'd0;
            rec_en                  <= 1'd0;
            rec_pkt_done            <= 1'd0;
        end
        else begin
            skip_en         <= 1'b0;
            error_en        <= 1'b0;
            rec_pkt_done    <= 1'b0;
            case(next_state)
                st_idle:begin
                    if((gmii_rx_dv == 1'b1) && (gmii_rxd == 8'h55))
                        skip_en <= 1'b1;        
                    else;
                end

                st_preamble:begin
                    if(gmii_rx_dv) begin
                        cnt <= cnt + 5'd1;
                        if((cnt < 5'd6) && (gmii_rxd != 8'h55))
                            error_en <= 1'b1;
                        else if(cnt == 5'd6) begin
                            cnt <= 5'd0;
                            if(gmii_rxd == 8'hd5) 
                                skip_en <= 1'b1;
                            else
                                error_en <= 1'b1;
                        end
                        else;
                    end
                    else;
                end

                st_eth_header:begin
                    if(gmii_rx_dv) begin
                        cnt <= cnt + 5'd1;
                        if(cnt < 5'd6)
                            des_mac <= {des_mac[39:0], gmii_rxd};
                        else if(cnt == 5'd12)
                            eth_type[15:8] <= gmii_rxd;
                        else if(cnt == 5'd13) begin
                            eth_type[7:0] <= gmii_rxd;
                            cnt <= 5'd0;
                            // �ж�MAC����̫������
                            if((des_mac == BOARD_MAC) || (des_mac == 48'hff_ff_ff_ff_ff_ff)
                            && (eth_type[15:8] == ETH_TYPE[15:8]) && (gmii_rxd == ETH_TYPE[7:0])) begin
                                skip_en <= 1'b1;
                            end
                            else
                                error_en <= 1'b1;
                        end
                        else;
                    end
                    else;
                end

                st_ip_header:begin
                    if(gmii_rx_dv) begin
                        cnt <= cnt + 5'd1;
                        if(cnt == 5'd0) 
                            ip_head_byte_num <= {gmii_rxd[3:0], 2'd0};              // IP�������ͷ�������ֶε�λ��4Bytes
                        else if(cnt == 5'd2) 
                            ip_total_length[15:8] <= gmii_rxd;
                        else if(cnt == 5'd3) 
                            ip_total_length[7:0]  <= gmii_rxd;                      
                        else if(cnt == 5'd4)
                            // ������Ч�����ֽڳ��ȣ�IPͷ20�ֽڣ�ICMPͷ8�ֽ�
                            icmp_data_length <= ip_total_length - 16'd28;
                        else if(cnt == 5'd9) begin
                            if(gmii_rxd != ICMP_TYPE) begin
                                error_en <= 1'b1;
                                cnt <= 5'd0;
                            end
                        end
                        else if((cnt >= 5'd16) && (cnt <= 5'd18))                  // ǰ�����ֽ�
                            des_ip <= {des_ip[23:0], gmii_rxd};
                        else if(cnt == 5'd19) begin
                            des_ip <= {des_ip[23:0], gmii_rxd};                    // ���һ���ֽ�
                            if((des_ip[23:0] == BOARD_IP[31:8]) && (gmii_rxd == BOARD_IP[7:0])) begin
                                skip_en <= 1'b1;
                                cnt <= 5'd0;
                            end
                            else begin
                                error_en <= 1'b1;
                                cnt <= 5'd0;
                            end
                        end
                        else;
                    end
                    else;
                end

                st_icmp_header:begin
                    if(gmii_rx_dv) begin
                        cnt <= cnt + 5'd1;
                        if(cnt == 5'd0)
                            icmp_type <= gmii_rxd;
                        else if(cnt == 5'd1)
                            icmp_code <= gmii_rxd;
                        else if(cnt == 5'd2) 
                            icmp_checksum[15:8] <= gmii_rxd;
                        else if(cnt == 5'd3)
                            icmp_checksum[7:0] <= gmii_rxd;
                        else if(cnt == 5'd4)
                            icmp_id[15:8] <= gmii_rxd;
                        else if(cnt == 5'd5)
                            icmp_id[7:0] <= gmii_rxd;
                        else if(cnt == 5'd6)
                            icmp_seq[15:8] <= gmii_rxd;
                        else if(cnt == 5'd7) begin
                            icmp_seq[7:0] <= gmii_rxd;
                            // �ж�ICMP�ı��������ǲ��ǻ�������
                            if(icmp_type  == ECHO_REQUEST) begin
                                skip_en <= 1'b1;
                                cnt <= 5'd0;
                            end
                            else begin
                                error_en <= 1'b1;                   // ICMP�������ʹ���
                                cnt <= 5'd0;
                            end
                        end
                        else;
                    end
                    else;
                end

                st_rx_data:begin
                    if(gmii_rx_dv) begin
                        rec_en_cnt <= rec_en_cnt + 2'd1;
                        icmp_rx_cnt <= icmp_rx_cnt + 16'd1;
                        rec_data <= gmii_rxd;
                        rec_en <= 1'b1;

                        // �жϽ��յ����ݸ�������ż������ÿ16bit����һ�μӷ�����
                        if(icmp_rx_cnt == icmp_data_length - 16'd1) begin
                            icmp_rx_data_d0 <= 8'h00;
                            if(icmp_data_length[0])
                                reply_checksum_add <= {8'd0, gmii_rxd} + reply_checksum_add;    // ���������
                            else
                                reply_checksum_add <= {icmp_rx_data_d0, gmii_rxd} + reply_checksum_add;     // �����ż��
                        end
                        else if(icmp_rx_cnt < icmp_data_length - 16'd1) begin           
                            icmp_rx_data_d0 <= gmii_rxd;
                            // icmp_rx_cnt <= icmp_rx_cnt + 16'd1;                        
                            if(icmp_rx_cnt[0] == 1'b1)
                                reply_checksum_add <= {icmp_rx_data_d0, gmii_rxd} + reply_checksum_add;
                            else
                                reply_checksum_add <= reply_checksum_add;
                        end
                        else;

                        if(icmp_rx_cnt == icmp_data_length - 16'd1) begin
                            skip_en <= 1'b1;
                            icmp_rx_cnt <= 16'd0;
                            rec_en_cnt <= 2'd0;
                            rec_pkt_done <= 1'b1;
                            rec_byte_num <= icmp_data_length;
                        end
                        else;
                    end
                    else;
                end

                st_rx_end:begin
                    rec_en <= 1'b0;
                    if(gmii_rx_dv == 1'b0 && skip_en == 1'b0) begin
                        reply_check_sum <= reply_checksum_add;
                        skip_en <= 1'b1;
                        reply_checksum_add <= 32'd0;
                    end
                    else;
                end
                
                default: ;
            endcase
        end
    end

endmodule
