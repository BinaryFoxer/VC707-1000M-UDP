`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// mdio����ģ��
//////////////////////////////////////////////////////////////////////////////////

module mdio_ctrl(
    input               clk,
    input               rst,

    input               soft_rst_trig,      // ��λ�����ź�
    input               op_done,            // ��������ź�
    input               op_rd_ack,          // ����Ӧ�ź�
    input       [15:0]  op_rd_data,         // �����ļĴ�������

    output  reg         op_exec,            // ��ʼ����
    output  reg         op_rh_wl,           // ��������
    output  reg [4:0]   op_addr,
    output  reg [15:0]  op_wr_data,         // д������

    output      [1:0]   led,                // �ٶ�ָʾled
    output              id_led,              // ��id��ȷָʾled
    output              test_led           // �����ʴ���ָʾled
    );

    // parameter define
    parameter READ_PERIOD = 24'd100_000;    // 20ms��һ��״̬�Ĵ���ֵ

    // reg define
    reg        rst_trig_0;
    reg        rst_trig_1;
    reg        rst_trig_2;
    reg        start_read;
    reg [23:0] timer_cnt;
    reg [4:0]  flow_cnt;
    reg [1:0]  speed_status;
    reg        rst_trig_flag;
    reg        link_error;
    reg [15:0] rd_data_t;
    reg [15:0] wr_data_t;
    reg        id_right;
    reg        test_led_v;

    // wire define
    wire pos_rst_trig;

    assign pos_rst_trig = ~rst_trig_2 & rst_trig_1;

    assign led = link_error ? 2'b00 : speed_status;
    assign id_led = id_right;
    // assign test_led = link_error;                         // ��PHY����ʧ��
    assign test_led = test_led_v;

    // ��soft_rst_trig�����ģ���ȡ������
    always @(posedge clk or posedge rst) begin
        if(rst)begin
            rst_trig_0 <= 0;
            rst_trig_1 <= 0;
            rst_trig_2 <= 0;
        end
        else begin
            rst_trig_0 <= soft_rst_trig;
            rst_trig_1 <= rst_trig_0;
            rst_trig_2 <= rst_trig_1;
        end
    end

    // ��ʱ��ȡ�ź�
    always @(posedge clk or posedge rst) begin
        if(rst)begin
            start_read <= 1'b0;
            timer_cnt <= 24'd0;
        end
        else begin
            if(timer_cnt == READ_PERIOD - 1) begin
                start_read <= 1'b1;
                timer_cnt <= 24'd0;
            end
            else begin
                timer_cnt <= timer_cnt + 24'd1;
                start_read <= 1'b0;
            end
        end
    end

    // ʹ�������������д���ƼĴ����Ͷ�״̬�Ĵ�������
    always @(posedge clk or posedge rst) begin
        if(rst)begin
            op_exec       <= 1'b0; 
            op_rh_wl      <= 1'b1;
            op_addr       <= 5'h0;
            op_wr_data    <= 16'd0;
            flow_cnt      <= 5'd0;
            speed_status  <= 2'b00;
            rst_trig_flag <= 1'b0;
            link_error    <= 1'b0;
            rd_data_t     <= 16'd0;
            wr_data_t     <= 16'd0;
            id_right      <= 1'b0;
            test_led_v    <= 1'b0;
        end
        else begin
            op_exec <= 1'b0;
            
            if(pos_rst_trig)
                rst_trig_flag <= 1'b1;
            case(flow_cnt)
                5'd0:begin
                    if(rst_trig_flag) begin                        // ʹ����λ����PHY���ã�д��Ĵ���
                        op_exec <= 1'b1;
                        op_rh_wl <= 1'b1;                          // ��R27����
                        op_addr <= 5'd27;                          // EPSSSR��ַ
                        flow_cnt <= 5'd1;       
                    end
                    else if(start_read) begin
                        op_exec <= 1'b1;
                        op_rh_wl <= 1'b1;                          // ������״̬�Ĵ���
                        op_addr <= 5'd1;                           // ����״̬�Ĵ���(BSCFR)��ַ
                        flow_cnt <= 5'd10;                         // �ȶ�phy id�����ԣ�
                        // test_led_v <= 1'b1;                        // ��ʼ��   
                    end                        
                end

                5'd1:begin
                    if(op_done) begin                              // �ȴ�R27���������
                        if(op_rd_ack == 1'b0) begin
                            rd_data_t <= op_rd_data;               // �Ĵ�R27��ʼ��������
                            flow_cnt <= 5'd2;                      
                        end
                        else
                            flow_cnt <= 5'd0;                      // R27���ʴ���
                                    
                    end
                end

                5'd2:begin
                    wr_data_t <= (rd_data_t & 16'b0111_1111_1111_0000) | 16'b1000_0000_0000_0000;   // ���ó�ǧ��SGMIIģʽ������λ����
                    flow_cnt <= 5'd3;
                end

                5'd3:begin
                    op_exec <= 1'b1;
                    op_rh_wl <= 1'b0;                              // дR27��������ģʽ
                    op_addr <= 5'd27;                              // EPSSSR��ַ
                    op_wr_data <= wr_data_t;                       // R27����������
                    flow_cnt <= 5'd4;
                end
                
                5'd4:begin
                    if(op_done) begin                              // �ȴ�дR27���
                        flow_cnt <= 5'd5;   
                    end
                end

                5'd5:begin
                    op_exec <= 1'b1;
                    op_rh_wl <= 1'b1;                        // �ȶ�R0�Ļ�������
                    op_addr <= 5'd0;
                    flow_cnt <= 5'd6;
                end

                5'd6:begin                                   
                    if(op_done) begin                       // �ȴ���R0���
                        if(op_rd_ack == 1'b0) begin
                            rd_data_t <= op_rd_data;
                            flow_cnt <= 5'd7;
                        end
                        else
                            flow_cnt <= 5'd0;               // R0���ʴ���
                                    
                    end
                end

                5'd7:begin
                    wr_data_t <= (rd_data_t & 16'b0000_0000_0011_1111) | 16'b1000_0001_0100_0000;       // bit[6]�����1Ϊ1000M����0Ϊ10M
                    flow_cnt <= 5'd8;
                end

                5'd8:begin
                    op_exec <= 1'b1;
                    op_rh_wl <= 1'b0;                          // ������ɣ���ʼд��λ
                    op_addr <= 5'd0;                           // �������ƼĴ���(BSCFR)��ַ
                    op_wr_data <= wr_data_t;     // ���ƼĴ�������: 1000_0001_0100_0000
                    flow_cnt <= 5'd9;
                end

                5'd9:begin
                    if(op_done) begin                           // ��λ��ɣ�������λ��־λ
                        flow_cnt <= 5'd0;
                        rst_trig_flag <= 1'b0;
                    end
                end

                // ------------��ʱ��״̬�Ĵ���-----------
                5'd10:begin
                    if(op_done) begin
                        if(op_rd_ack == 1'b0 && op_rd_data[2] == 1) begin  // ����Ӧ�Լ��������� && op_rd_data[2] == 1��op_rd_ack == 1'b0
                            flow_cnt <= 5'd11;
                            link_error <= 1'b0;
                            test_led_v <= 1'b1;
                        end
                        else begin
                            flow_cnt <= 5'd0;
                            link_error <= 1'b1;
                        end
                    end
                    else begin
                        // link_error <= 1'b1;                               // ���û�ж���Ӧ��Ҳ��������ʧ��(����)
                        // test_led_v <= 1'b1;
                    end
                end

                5'd11:begin
                    op_exec <= 1'b1;
                    op_rh_wl <= 1'b1;                        // ��PHY״̬�Ĵ���
                    op_addr <= 5'd17;                        // PHY״̬�Ĵ���R17��ַ
                    flow_cnt <= 5'd12;
                end

                5'd12:begin
                    if(op_done) begin
                        if(op_rd_ack == 1'b0)                // �ж���Ӧ��˵�����ɹ���������
                            flow_cnt <= 5'd13;
                        else
                            flow_cnt <= 5'd0;
                    end
                end

                5'd13:begin
                    case(op_rd_data[15:14])
                        2'b00:speed_status <= 2'b01;    // 10mbps
                        2'b01:speed_status <= 2'b10;    // 100mbps
                        2'b10:speed_status <= 2'b11;    // 1000mbps
                        default:speed_status <= 2'b00;
                    endcase
                    flow_cnt <= 5'd14;                   
                end

                5'd14:begin
                    op_exec <= 1'b1;                        // �����phy ID״̬��ȷ����������оƬ����
                    op_rh_wl <= 1'b1;                       // ��PHY ID�Ĵ���
                    op_addr <= 5'd2;                        // �Ĵ���R2��ַ
                    flow_cnt <= 5'd15;
                end

                5'd15:begin
                    if(op_done) begin
                        if(op_rd_ack == 1'b0) begin
                            rd_data_t <= op_rd_data;
                            flow_cnt <= 5'd16;
                        end
                        else
                            flow_cnt <= 5'd0;
                    end
                end

                5'd16:begin
                    flow_cnt <= 5'd0;
                    id_right <= (rd_data_t == 16'h0141) ? 1'b1 : 1'b0;
                    // test_led_v <= 1'b1;
                end

            endcase
        end
    end


endmodule
