`timescale 1ns / 1ps

// ----------------------------------------------------------------
// ���գ����Զ˷�������gmii_rxd
// ���ܣ����mac֡�Ľ��գ�����mac֡�ṹ�жϽ����Ƿ���ȷ/�Ƿ�ΪĿ�ķ�
// ���CRC32���У��
// ----------------------------------------------------------------

module arp_rx(
    input                   rst,            // ϵͳ��λ                
    input                   clk,            // ������gmii����ʱ��
    
    input                   gmii_rx_dv,     // gmii����������Ч
    input          [7:0]    gmii_rxd,       // gmii��������

    output reg              arp_rx_done,    // arp�������ݴ������
    output reg              arp_rx_type,    // arp�����������ͣ�����/Ӧ��
    output reg     [31:0]   src_ip,         // ���ͷ�Դip��ַ
    output reg     [47:0]   src_mac,        // ���ͷ�Դmac��ַ
    output reg              arp_get,
    output reg     [4:0]    cur_state
    );

    // parameter define
    parameter  BOARD_MAC = 48'h00_11_22_33_44_55;        // �忨MAC��ַ
    parameter  BOARD_IP  = {8'd192,8'd168,8'd0,8'd2};
    
    localparam ETH_TYPE     = 16'h08_06;                    // ��̫��֡���͡�ARP֡Ϊ0806
    localparam st_idle      = 5'b0_0001;
    localparam st_preamble  = 5'b0_0010;
    localparam st_header    = 5'b0_0100;
    localparam st_arp_data  = 5'b0_1000;
    localparam st_arp_end   = 5'b1_0000;

    // reg define
    // reg [4:0]   cur_state;
    reg [4:0]   next_state;
    reg [4:0]   cnt;                      // �������յ��ֽ�
    reg         skip_en;                  // ״̬��תʹ��
    reg         error_en;                 // ������תʹ��
    reg [47:0]  des_mac_t;                // �Ĵ���յ���Ŀ��mac
    reg [31:0]  des_ip_t;                 // �Ĵ���յ���Ŀ��ip
    reg [15:0]  eth_type_t;               // �Ĵ���յ�����̫֡����
    reg [15:0]  op_code;                  // ������
    reg [47:0]  src_mac_t;                // �Ĵ���յ���Դmac
    reg [31:0]  src_ip_t;                 // �Ĵ���յ���Դip 
    reg         rx_done_t;                // �Ĵ�arp�������ݴ�������ź�                             


    // ----------------------------arp����֡����----------------------------
    // ͬ��ʱ������״̬ת��
    always @(posedge clk or posedge rst) begin
        if(rst) 
            cur_state <= st_idle;
        else
            cur_state <= next_state;
    end

    // ����߼�����״̬ת������
    always @(*) begin
        next_state = cur_state;
        case (cur_state)
            st_idle:begin
                if(skip_en) 
                    next_state = st_preamble;
                else
                    next_state = st_idle;
            end

            st_preamble:begin
                if(skip_en)
                    next_state = st_header;
                else if(error_en)
                    next_state = st_arp_end;
                else
                    next_state = st_preamble;
            end

            st_header:begin
                if(skip_en)
                    next_state = st_arp_data;
                else if(error_en)
                    next_state = st_arp_end;
                else
                    next_state = st_header;
            end

            st_arp_data:begin
                if(skip_en)
                    next_state = st_arp_end;
                else if(error_en)
                    next_state = st_arp_end;
                else   
                    next_state = st_arp_data;
            end

            st_arp_end:begin
                if(skip_en)
                    next_state = st_idle;
                else
                    next_state = st_arp_end;
            end

            default: next_state = st_idle;
        endcase
    end

    // ͬ��ʱ������״̬���
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            cnt         <= 5'd0;
            skip_en     <= 1'd0;
            error_en    <= 1'd0;
            des_mac_t   <= 48'd0;
            des_ip_t    <= 32'd0;
            eth_type_t  <= 16'd0;
            op_code     <= 16'd0;
            src_mac_t   <= 48'd0;
            src_ip_t    <= 32'd0;
            rx_done_t   <= 1'd0;
            arp_rx_type <= 1'd0;
            src_ip      <= 32'd0;
            src_mac     <= 48'd0;
            arp_get     <= 1'b0;
        end
        else begin
            skip_en <= 1'b0;
            error_en <= 1'b0;
            rx_done_t <= 1'b0;
            arp_get   <= 1'b0;
            case(next_state)                                        // ��Ҫcur_state��ת������������������next_state
                st_idle:begin
                    if((gmii_rx_dv == 1) && (gmii_rxd == 8'h55)) begin
                        skip_en <= 1'b1;                            // ����������Ч���Ҽ�⵽ǰ����
                    end
                end

                st_preamble:begin
                    if(gmii_rx_dv == 1'b1) begin
                        cnt <= cnt + 5'd1;
                        if((cnt < 5'd6) && (gmii_rxd != 8'h55)) 
                            error_en <= 1'b1;               // ���ǰ�߸��ֽ����Ѿ����ִ���
                        else if(cnt == 5'd6) begin
                            cnt <= 5'b0;
                            if(gmii_rxd == 8'hd5)begin           // �ڰ˸��ֽڼ�⵽��ʼ�ַ�
                                skip_en <= 1'b1;
                            end
                            else
                                error_en <= 1'b1;
                        end
                    end
                end

                st_header:begin                            // �ж�Ŀ��mac��֡����
                    if(gmii_rx_dv == 1'b1) begin
                        cnt <= cnt + 5'd1;
                        if(cnt < 5'd6) 
                            des_mac_t <= {des_mac_t[39:0], gmii_rxd};   // ����Ŀ��mac
                        else if(cnt == 5'd6) begin
                            if((des_mac_t != BOARD_MAC) && des_mac_t != 48'hff_ff_ff_ff_ff_ff)           
                                error_en <= 1'b1;         // Ŀ��mac���ǰ忨���Ҳ��ǹ㲥��ַ  
                        end
                        else if(cnt == 5'd12) 
                            eth_type_t[15:8] <= gmii_rxd;  // ����֡����
                        else if(cnt == 5'd13) begin
                            cnt <= 5'd0;
                            eth_type_t[7:0] <= gmii_rxd;   // ����֡����
                            if((eth_type_t[15:8] == ETH_TYPE[15:8]) && 
                                (gmii_rxd == ETH_TYPE[7:0])) begin
                                    skip_en <= 1'b1;
                                    
                                end            // �ж��Ƿ���ARP���� 
                            else
                                error_en <= 1'b1;
                        end
                    end
                end

                st_arp_data:begin
                    if(gmii_rx_dv == 1'b1) begin
                        cnt <= cnt + 5'd1;
                        if(cnt == 5'd6)                                 // ������
                            op_code[15:8] <= gmii_rxd;
                        else if(cnt == 5'd7)
                            op_code[7:0] <= gmii_rxd;
                        else if(cnt >= 5'd8 && cnt < 5'd14)             // Դmac
                            src_mac_t <= {src_mac_t[39:0], gmii_rxd};
                        else if(cnt >= 5'd14 && cnt < 5'd18)            // Դip
                            src_ip_t <= {src_ip_t[23:0], gmii_rxd};
                        else if(cnt >= 5'd24 && cnt < 5'd28)            // Ŀ��ip
                            des_ip_t <= {des_ip_t[23:0], gmii_rxd};
                        else if(cnt == 5'd28) begin
                            cnt <= 5'd0;
                            if(des_ip_t == BOARD_IP) begin
                                arp_get <= 1'b1;
                                if(op_code == 16'd1 || op_code == 16'd2) begin
                                    skip_en   <= 1'b1;
                                    rx_done_t <= 1'b1;
                                    src_mac   <= src_mac_t;
                                    src_ip    <= src_ip_t;
                                    src_mac_t <= 48'd0;
                                    src_ip_t  <= 32'd0;
                                    des_mac_t <= 48'd0;
                                    des_ip_t  <= 32'd0;
                                    if(op_code == 16'd1)
                                        arp_rx_type <= 1'b0;            // arp����
                                    else
                                        arp_rx_type <= 1'b1;            // arpӦ��
                                end
                                else
                                    error_en <= 1'b1;
                            end
                            else  
                                error_en <= 1'b1;
                        end
                    end
                end

                st_arp_end:begin
                    cnt <= 5'd0;
                    // ���������ݽ������
                    if(gmii_rx_dv == 1'b0 && skip_en == 1'b0)
                        skip_en <= 1'b1;    
                end
            default: ;
            endcase
        end
    end

// ���arp_rx_done�ź�
always @(posedge clk or posedge rst) begin
    if(rst)
        arp_rx_done <= 1'b0;
    else
        arp_rx_done <= rx_done_t;
end

endmodule
