`timescale 1ns / 1ps

// --------------------------------------------------------------------
// UDP��������ģ��
// ��ǰ����UDP���ز���
// --------------------------------------------------------------------

module eth_udp_test(
    input               sys_clk_p,               // 200mhzʱ��Դ
    input               sys_clk_n,
    input               sys_rst,

    // --------mdio�ӿ�--------
    output              eth_mdc,
    inout               eth_mdio,

    output      [1:0]   led,
    output              id_led,              // ��id��ȷָʾled
    output              test_led,            // �����ʴ���ָʾled
    output              download_sus,        // ���ش���ɹ�ָʾled
    input               touch_key,           // mdio���ð���

    // --------SGMII�ӿ�-------
    input               sgmii_clk_n,             // 125m�ο�ʱ��
    input               sgmii_clk_p,
    input               sgmii_rxn,                      
    input               sgmii_rxp,
    output              sgmii_txn,
    output              sgmii_txp,              
    output              eth_rst_n,               // ��̫��ģ�鸴λ

    input               send_key,                // ����arp���󰴼�
    output              arp_led                  // arp����led

    );

    // �忨mac��ip
    parameter  BOARD_MAC = 48'h00_11_22_33_44_55;        // �忨MAC��ַ
    parameter  BOARD_IP  = {8'd192,8'd168,8'd0,8'd2}; 
    // Ŀ��mac��ip
    parameter  DES_MAC   = 48'hff_ff_ff_ff_ff_ff;
    parameter  DES_IP  = {8'd192,8'd168,8'd0,8'd3}; 

    // wire define
    wire                gmii_tx_en;
    wire                gmii_tx_er;
    wire        [7:0]   gmii_txd;
    wire                gmii_tx_clk;
    wire                gmii_tx_done;
    wire                gmii_rx_clk;
    wire                gmii_rx_dv;
    wire                gmii_rx_er;
    wire        [7:0]   gmii_rxd;

    wire                arp_gmii_tx_en;
    wire        [7:0]   arp_gmii_txd;
    wire                arp_tx_en;
    wire                arp_tx_type;
    wire                arp_tx_done;
    wire                arp_rx_done;
    wire                arp_rx_type;

    wire                resetdone;
    wire                mmcm_locked_out;
    wire        [47:0]  des_mac;
    wire        [31:0]  des_ip;
    wire        [31:0]  src_ip;
    wire        [47:0]  src_mac;
    wire                sys_clk;

    wire                sgmii_clk_en;
    wire        [15:0]  status_vector;
    wire                arp_get;
    wire        [4:0]   cur_state;  

    // ICMP�˿��ź�
    wire                icmp_tx_start_en;              // ICMP����ģ��ʹ���źţ���ʼ�����
    wire                icmp_tx_done;                  // ICMP�����������
    wire                icmp_gmii_tx_en;               // ICMPʹ��gmii_txd��������
    wire        [7:0]   icmp_gmii_txd;                 // ICMPͨ��gmii_txd���͵�����
    wire                icmp_rec_en;                   // ICMP��������ʹ���ź�
    wire        [7:0]   icmp_rec_data;
    wire                icmp_tx_req;                   // ICMP�����������ź�
    wire        [7:0]   icmp_tx_data;                  // ICMP����������
    wire                icmp_rec_pkt_done;
    wire        [15:0]  icmp_rec_byte_num;             // ������Ч�ֽ���     
    wire        [15:0]  icmp_tx_byte_num;              // ������Ч�ֽ���

    // UDP�˿��ź�
    wire                udp_gmii_tx_en;
    wire        [7:0]   udp_gmii_txd;

    wire                udp_rec_pkt_done;              // �������ݰ���ɱ�־
    wire                udp_rec_en;                    // ��������ʹ��
    wire        [7:0]   udp_rec_data;                  // udp��������
    wire        [15:0]  udp_rec_byte_num;              // ������Ч�ֽ���
    wire                udp_tx_start_en;               // ��ʼ���ʹ����ź�
    wire        [7:0]   udp_tx_data;                   // udp��������        
    wire        [15:0]  udp_tx_byte_num;               // ������Ч�ֽ���
    wire                udp_tx_done;                   // ��������ź�
    wire                udp_tx_req;                    // ��ȡ�������������ź�

    wire        [7:0]   rec_data;
    wire                rec_en;
    wire        [7:0]   tx_data;
    wire                tx_req;

    assign  icmp_tx_start_en = icmp_rec_pkt_done;
    assign  icmp_tx_byte_num = icmp_rec_byte_num;

    assign  udp_tx_start_en = udp_rec_pkt_done;
    assign  udp_tx_byte_num = udp_rec_byte_num;
    assign  des_ip = src_ip;
    assign  des_mac = src_mac;
    assign  eth_rst_n = ~sys_rst;

    assign download_sus = arp_get;

    // ----------------------   ila����   ------------------------
    ila_1 icmp_ila_test_1 (
        .clk(gmii_tx_clk), // input wire clk
    
        .probe0(icmp_tx_start_en), // input wire [0:0]  probe0  
        .probe1(tx_req), // input wire [0:0]  probe1 
        .probe2(rec_en), // input wire [0:0]  probe2 
        .probe3(gmii_rx_dv), // input wire [0:0]  probe3 
        .probe4(gmii_rxd), // input wire [7:0]  probe4 
        .probe5(gmii_txd), // input wire [7:0]  probe5 
        .probe6(icmp_gmii_txd), // input wire [7:0]  probe6 
        .probe7(icmp_rec_byte_num), // input wire [15:0]  probe7 
        .probe8(icmp_tx_done), // input wire [0:0]  probe8 
        .probe9(udp_tx_done), // input wire [0:0]  probe9 
        .probe10(rec_data), // input wire [7:0]  probe10 
        .probe11(tx_data), // input wire [7:0]  probe11
        .probe12(cur_state)
    );

    // ---------------------------------����200mhzʱ��Դ-------------------------------------
    IBUFDS #(
      .DIFF_TERM("FALSE"),       // Differential Termination
      .IBUF_LOW_PWR("FALSE"),     // Low power="TRUE", Highest performance="FALSE" 
      .IOSTANDARD("LVDS")     // Specify the input I/O standard
   ) IBUFDS_inst (
      .O(sys_clk),  // Buffer output
      .I(sys_clk_p),  // Diff_p buffer input (connect directly to top-level port)
      .IB(sys_clk_n) // Diff_n buffer input (connect directly to top-level port)
   );

    // arpģ������
    arp #(
        .DES_IP             (DES_IP),
        .DES_MAC            (DES_MAC),
        .BOARD_IP           (BOARD_IP),
        .BOARD_MAC          (BOARD_MAC)
    )u_arp(
        .rst                (sys_rst),          
        .gmii_rx_clk        (gmii_tx_clk),
        .gmii_rx_dv         (gmii_rx_dv), 
        .gmii_rxd           (gmii_rxd),   
        .gmii_tx_clk        (gmii_tx_clk),
        .gmii_tx_en         (arp_gmii_tx_en), 
        .gmii_txd           (arp_gmii_txd),   
        .gmii_tx_done       (arp_tx_done),              

        .arp_tx_en          (arp_tx_en),  
        .arp_tx_type        (arp_tx_type),
        .arp_rx_done        (arp_rx_done),
        .arp_rx_type        (arp_rx_type),
        .des_mac            (des_mac),    
        .des_ip             (des_ip),     
        .src_mac            (src_mac),    
        .src_ip             (src_ip),
        
        .arp_led            (arp_led),
        .arp_get            (arp_get),
        .cur_state          (cur_state)  
    );

    // ICMPģ������
    icmp #(
        .BOARD_IP(BOARD_IP),
        .BOARD_MAC(BOARD_MAC),
        .DES_IP(DES_IP),
        .DES_MAC(DES_MAC)
    )u_icmp(
        .rst                (sys_rst        ),
        .gmii_rx_clk        (gmii_tx_clk    ),
        .gmii_rx_dv         (gmii_rx_dv     ),
        .gmii_rxd           (gmii_rxd       ),
        .gmii_tx_clk        (gmii_tx_clk    ),
        .gmii_tx_en         (icmp_gmii_tx_en),
        .gmii_txd           (icmp_gmii_txd  ),
        .rec_pkt_done       (icmp_rec_pkt_done),
        .rec_en             (icmp_rec_en    ),
        .rec_data           (icmp_rec_data  ),
        .rec_byte_num       (icmp_rec_byte_num),
        .tx_start_en        (icmp_tx_start_en),
        .tx_data            (icmp_tx_data   ),
        .tx_byte_num        (icmp_tx_byte_num),
        .des_mac            (des_mac        ),
        .des_ip             (des_ip         ),
        .tx_done            (icmp_tx_done   ),
        .tx_req             (icmp_tx_req    )
    );

    // ͬ��FIFO����
    fifo_generator_0 data_fifo (
      .clk(gmii_tx_clk),      // input wire clk
      .srst(sys_rst),    // input wire srst
      .din(rec_data),      // input wire [7 : 0] din
      .wr_en(rec_en),  // input wire wr_en
      .rd_en(tx_req),  // input wire rd_en
      .dout(tx_data),    // output wire [7 : 0] dout
      .full(),    // output wire full
      .empty()  // output wire empty
    );

    eth_ctrl_sw u_eth_ctrl_sw(
        .clk                (gmii_tx_clk),
        .rst                (sys_rst),

        // ARP�˿��ź�
        .arp_rx_done        (arp_rx_done),                   // ARP���ݰ���������ź�
        .arp_rx_type        (arp_rx_type),                   // ARP�������ͣ�0������1��Ӧ��
        .arp_tx_en          (arp_tx_en),                     // ARP����ģ��ʹ���źţ���ʼ�����
        .arp_tx_type        (arp_tx_type),                   // ARP�������ͣ�0������1��Ӧ��
        .arp_tx_done        (arp_tx_done),                   // ARP�����������
        .arp_gmii_tx_en     (arp_gmii_tx_en),                // ARPʹ��gmii_txd��������
        .arp_gmii_txd       (arp_gmii_txd),                  // ARPͨ��gmii_txd���͵�����

        // ICMP�˿��ź�
        .icmp_tx_start_en   (icmp_tx_start_en),              // ICMP����ģ��ʹ���źţ���ʼ�����
        .icmp_tx_done       (icmp_tx_done),                  // ICMP�����������
        .icmp_gmii_tx_en    (icmp_gmii_tx_en),               // ICMPʹ��gmii_txd��������
        .icmp_gmii_txd      (icmp_gmii_txd),                 // ICMPͨ��gmii_txd���͵�����

        // ICMP fifo�ӿ��ź�
        .icmp_rec_en        (icmp_rec_en),                   // ICMP��������ʹ���ź�
        .icmp_rec_data      (icmp_rec_data),
        .icmp_tx_req        (icmp_tx_req),                   // ICMP�����������ź�
        .icmp_tx_data       (icmp_tx_data),                  // ICMP����������

        // UDP��ض˿��ź�
        .udp_tx_start_en    (udp_tx_start_en),               // UDP����ģ��ʹ���źţ���ʼ�����
        .udp_tx_done        (udp_tx_done),                   // UDP��������ź�
        .udp_gmii_tx_en     (udp_gmii_tx_en),                // UDPʹ��gmii_txd��������
        .udp_gmii_txd       (udp_gmii_txd),                  // UDPͨ��gmii_txd���͵�����

        // UDP fifo�ӿ��ź�
        .udp_rec_en         (udp_rec_en),                   // UDP��������ʹ���ź�
        .udp_rec_data       (udp_rec_data),
        .udp_tx_req         (udp_tx_req),                   // UDP�����������ź�
        .udp_tx_data        (udp_tx_data),                  // UDP����������

        // fifo�ӿ��ź�
        .tx_data            (tx_data),                      // ����������
        .tx_req             (tx_req),
        .rec_en             (rec_en),
        .rec_data           (rec_data),

        // GMII��������
        .gmii_tx_en         (gmii_tx_en),
        .gmii_txd           (gmii_txd)
    );

    udp #(
        .BOARD_IP(BOARD_IP),
        .BOARD_MAC(BOARD_MAC),
        .DES_IP(DES_IP),
        .DES_MAC(DES_MAC)
    )u_udp(
        .rst                    (sys_rst),
        // GMII�ӿ�
        .gmii_rx_clk            (gmii_tx_clk),
        .gmii_rx_dv             (gmii_rx_dv),
        .gmii_rxd               (gmii_rxd),
        .gmii_tx_clk            (gmii_tx_clk),
        .gmii_tx_en             (udp_gmii_tx_en),
        .gmii_txd               (udp_gmii_txd),

        // �û��ӿ�
        .rec_pkt_done           (udp_rec_pkt_done),               // �������ݰ���ɱ�־
        .rec_en                 (udp_rec_en),                     // ��������ʹ��
        .rec_data               (udp_rec_data),                   // udp��������
        .rec_byte_num           (udp_rec_byte_num),               // ������Ч�ֽ���
        .tx_start_en            (udp_tx_start_en),                // ��ʼ���ʹ����ź�
        .tx_data                (udp_tx_data),                    // udp��������        
        .tx_byte_num            (udp_tx_byte_num),                // ������Ч�ֽ���
        .des_mac                (des_mac),
        .des_ip                 (des_ip),
        .tx_done                (udp_tx_done),                    // ��������ź�
        .tx_req                 (udp_tx_req)                      // ��ȡ�������������ź�

    );

    // sgmii gmii�ӿ�ת������
    sgmii_to_gmii u_sgmii_gmii(
        .sys_rst                    (sys_rst    ),             
        .sgmii_clk_n                (sgmii_clk_n),   
        .sgmii_clk_p                (sgmii_clk_p),   
        .independent_clock_bufg     (sys_clk    ),
        .sgmii_rx_n                 (sgmii_rxn  ),    
        .sgmii_rx_p                 (sgmii_rxp  ),    
        .gmii_tx_en                 (gmii_tx_en ),    
        .gmii_tx_er                 (),    
        .gmii_txd                   (gmii_txd   ),                            
        .gmii_rx_clk                (gmii_rx_clk),   
        .gmii_rx_dv                 (gmii_rx_dv ),    
        .gmii_rx_er                 (),    
        .gmii_rxd                   (gmii_rxd   ),      
        .gmii_tx_clk                (gmii_tx_clk),   
        .sgmii_tx_n                 (sgmii_txn  ),    
        .sgmii_tx_p                 (sgmii_txp  ),                          
        .resetdone                  (resetdone  ),     
        .mmcm_locked_out            (mmcm_locked_out),
        .sgmii_clk_en               (sgmii_clk_en),
        .status_vector              (status_vector)

    );

    // mdio����ӿ�����
    mdio_wr_test u_mdio_wr_test(
        .sys_clk(sys_clk),
        .sys_rst(sys_rst),
        .eth_rst_n(eth_rst_n),
        .eth_mdc(eth_mdc),
        .eth_mdio(eth_mdio),
        .touch_key(touch_key),
        .led(led),
        .id_led(id_led),
        .test_led(test_led)
    );



endmodule
