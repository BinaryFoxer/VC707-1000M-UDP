`timescale 1ns / 1ps

module mac_send(
    // �����ź�
    input tx_go,
    input rst_n,
    input [10:0] pyd_length,   //payload�������ݳ���
    
    // mac֡ͷ
    input [47:0] src_mac,
    input [47:0] des_mac,
    input [15:0] type_length,
    
    // mac�����غ�
    output reg fifo_rdreq,
    input [7:0] fifo_rddata,
    input fifo_rdclk,
    
    // CRCУ����
    input [31:0] crc_result,
    
    // gmii���ݴ���ӿ�
    input gmii_clk,
    output reg gmii_tx_en,
    output reg gmii_tx_err,
    output reg [7:0] gmii_tx_data
    
    );
    
    // ====================�Ĵ������==================
    reg [5:0] cnt;  // �����ֽڼ����߼�
    reg en_cnt; // ״̬����ʹ���źţ�������23��ȡFIFOʱ�ü���ֹͣ����
    reg [10:0] pyd_data_num;    // payload�ֽڼ���
    reg en_tx;
    
    parameter CRC32 = 32'h967D1D69;
    assign crc_result = {CRC32[7:0], CRC32[15:8], CRC32[23:16], CRC32[31:24]};
    
    // =================���л������߼�==================
    always@(posedge gmii_clk or negedge rst_n) begin
        if(!rst_n) begin
            gmii_tx_data <= 8'd0;
        end else begin
            case(cnt)
                1, 2, 3, 4, 5, 6, 7:
                     gmii_tx_data <= 8'h55;     // ǰ����
                     
                8: gmii_tx_data <= 8'hd5;       // �ָ���
                // Ŀ��mac
                9: gmii_tx_data <= des_mac[47:40];
                10: gmii_tx_data <= des_mac[39:32];
                11: gmii_tx_data <= des_mac[31:24];
                12: gmii_tx_data <= des_mac[23:16];
                13: gmii_tx_data <= des_mac[15:8];
                14: gmii_tx_data <= des_mac[7:0];
                // Դmac
                15: gmii_tx_data <= src_mac[47:40];
                16: gmii_tx_data <= src_mac[39:32];
                17: gmii_tx_data <= src_mac[31:24];
                18: gmii_tx_data <= src_mac[23:16];
                19: gmii_tx_data <= src_mac[15:8];
                20: gmii_tx_data <= src_mac[7:0];
                // ���ͳ���
                21: gmii_tx_data <= type_length[15:8];
                22: gmii_tx_data <= type_length[7:0];
                // ��fifo�ж�ȡpayload
                23: gmii_tx_data <= fifo_rddata;
                
                24: gmii_tx_data <= crc_result[31:24];
                25: gmii_tx_data <= crc_result[23:16];
                26: gmii_tx_data <= crc_result[15:8];
                27: gmii_tx_data <= crc_result[7:0];
                
                // ����֡����
                28: gmii_tx_data <= 8'd0;
                default: gmii_tx_data <= 8'd0;
         
            endcase
        
        end
        
    end
    
    // ================����ֵ23ʱ��FIFO��������==============
    // en_cntû����ʱһ�ģ����̾�������
    assign en_cnt = !((cnt==23) && (pyd_data_num>1));  //����ֹͣ����ȡfifo���ݵ�����
    assign fifo_rdreq = !en_cnt;
    
//    // fifo_rdreq����һ��
//    always@(posedge gmii_clk or negedge rst_n) begin
//        if(!rst_n) begin
//            fifo_rdreq <= 1'd0;     
//        end else if(!en_cnt) begin
//                fifo_rdreq <= 1'd1;   
//        end else begin
//            fifo_rdreq <= 1'd0;
//        end
        
//    end
    
    // �ö�ȡ���ݳ��ȿ��ƶ�ȡfifoʱ��
    always@(posedge gmii_clk or negedge rst_n) begin
        if(!rst_n) begin
            pyd_data_num <= 11'd0;
        end else if(tx_go) begin    // tx_go��һ�������źţ�ֻ�ڿ�ʼ����ʱ���1�θߵ�ƽ
            pyd_data_num <= pyd_length;      
        end else if(!en_cnt) begin
                pyd_data_num <= pyd_data_num - 11'd1;   
        end else begin
            pyd_data_num <= pyd_data_num;
        end
     
    end
    
    // =================cnt�����߼�==================
    // �ڲ�����ʹ�ܣ�ʵ�ʷ���ʱ�䲻���з��ͼ����ô��
    always@(posedge gmii_clk or negedge rst_n) begin
        if(!rst_n)
            en_tx <= 1'b0;
        else if(tx_go) 
            en_tx <= 1'b1;
        else if(cnt >= 6'd27)
            en_tx <= 1'b0;
        else 
            en_tx <= en_tx;
       
    end
    
    always@(posedge gmii_clk or negedge rst_n) begin
        if(!rst_n)
            cnt <= 5'd0;
        else if(en_tx) begin
            if(!en_cnt) 
                cnt <= cnt;
            else 
                cnt <= cnt + 6'd1;
        end else begin
            cnt <= 6'd0;
        end
    
    end
    
    // =====================gmiiתsgmii���ٴ��нӿ�========================
    // VC707�������֧��sgmii�ӿڴ���
    

    
    
   
endmodule



