`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// mdio����ģ��
//////////////////////////////////////////////////////////////////////////////////

module soft_rst_only(
    input               clk,
    input               rst_n,

    input               soft_rst_trig,      // ��λ�����ź�
    input               op_done,            // ��������ź�
    input               op_rd_ack,          // ����Ӧ�ź�
    input       [15:0]  op_rd_data,         // �����ļĴ�������

    output  reg         op_exec,            // ��ʼ����
    output  reg         op_rh_wl,           // ��������
    output  reg [4:0]   op_addr,
    output  reg [15:0]  op_wr_data,         // д������

    output      [1:0]   led                 // �ٶ�ָʾled
    );

    // parameter define
    parameter READ_PERIOD = 24'd100_000;    // 10ms��һ��״̬�Ĵ���ֵ

    // reg define
    reg        rst_trig_0;
    reg        rst_trig_1;
    reg        rst_trig_2;
    reg        start_read;
    reg [23:0] timer_cnt;
    reg [3:0]  flow_cnt;
    reg [1:0]  speed_status;
    reg        rst_trig_flag;
    reg        link_error;

    // wire define
    wire pos_rst_trig;

    assign pos_rst_trig = ~rst_trig_2 & rst_trig_1;

    assign led = link_error ? 2'b00 : speed_status;

    // ��soft_rst_trig�����ģ���ȡ������
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n)begin
            rst_trig_0 <= 0;
            rst_trig_1 <= 0;
            rst_trig_2 <= 0;
        end
        else begin
            rst_trig_0 <= soft_rst_trig;
            rst_trig_1 <= rst_trig_0;
            rst_trig_2 <= rst_trig_1;
        end
    end

    // ��ʱ��ȡ�ź�
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n)begin
            start_read <= 1'b0;
            timer_cnt <= 24'd0;
        end
        else begin
            if(timer_cnt == READ_PERIOD - 1) begin
                start_read <= 1'b1;
                timer_cnt <= 24'd0;
            end
            else begin
                timer_cnt <= timer_cnt + 24'd1;
                start_read <= 1'b0;
            end
        end
    end

    // ʹ�������������д���ƼĴ����Ͷ�״̬�Ĵ�������
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n)begin
            op_exec       <= 1'b0; 
            op_rh_wl      <= 1'b1;
            op_addr       <= 5'h0;
            op_wr_data    <= 16'd0;
            flow_cnt      <= 4'd0;
            speed_status  <= 2'b00;
            rst_trig_flag <= 1'b0;
            link_error    <= 1'b0;
        end
        else begin
            op_exec <= 1'b0;
            if(pos_rst_trig)
                rst_trig_flag <= 1'b1;
            case(flow_cnt)
                4'd0:begin
                    if(rst_trig_flag) begin
                        op_exec <= 1'b1;
                        op_rh_wl <= 1'b0;                          // д��λ
                        op_addr <= 5'd0;                           // �������ƼĴ���(BSCFR)��ַ
                        op_wr_data <= 16'b1010_0001_0100_0000;     // ���ƼĴ�������: 1010_0001_0100_0000
                        flow_cnt <= 4'd1;       
                    end
                    else if(start_read) begin
                        op_exec <= 1'b1;
                        op_rh_wl <= 1'b1;                          // ������״̬�Ĵ���
                        op_addr <= 5'd1;                           // ����״̬�Ĵ���(BSCFR)��ַ
                        flow_cnt <= 4'd2;   
                    end                        
                end

                4'd1:begin
                    if(op_done)                             // ��λ��ɣ�������λ��־λ
                        flow_cnt <= 4'd0;
                        rst_trig_flag <= 4'd0;
                end

                4'd2:begin
                    if(op_done) begin
                        if(op_rd_ack == 1'b0 && op_rd_data[5] == 1'b1 && op_rd_data[2] == 1'b1) begin  // ����Ӧ����Э���Լ���������
                            flow_cnt <= 4'd3;
                            link_error <= 1'b0;
                        end
                        else begin
                            flow_cnt <= 4'd0;
                            link_error <= 1'b1;
                        end
                    end
                end

                4'd3:begin
                    op_exec <= 1'b1;
                    op_rh_wl <= 1'b1;                        // ��PHY״̬�Ĵ���
                    op_addr <= 5'd2;                        // PHY״̬�Ĵ���R17��ַ�����Զ�phy_id1
                    flow_cnt <= 4'd4;
                end

                4'd4:begin
                    if(op_done) begin
                        if(op_rd_ack == 1'b0)                // �ж���Ӧ��˵�����ɹ���������
                            flow_cnt <= 4'd5;
                        else
                            flow_cnt <= 4'd0;
                    end
                end

                4'd5:begin
                    flow_cnt <= 4'd0;
                    case(op_rd_data[15:14])
                        2'b00:speed_status <= 2'b01;    // 10mbps
                        2'b01:speed_status <= 2'b10;    // 100mbps
                        2'b10:speed_status <= 2'b11;    // 1000mbps
                        default:speed_status <= 2'b00;
                    endcase
                end
            endcase
        end
    end



endmodule
