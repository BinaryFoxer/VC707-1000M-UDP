`timescale 1ns / 1ps

module arp_send(
    input rst_n,
    input gmii_clk,
    
    // gmii�ӿ�
    output reg gmii_tx_err,
    output reg gmii_tx_en,
    output reg [7:0] gmii_tx_data

    );
    
    // ============���������=================
    reg [24:0] cnt;

    
    // ===========mac_sendʵ����================
        // �����ź�
    wire tx_go;
    // mac�����غ�
    reg fifo_rdreq;
    reg [7:0] fifo_rddata;
    reg fifo_rdclk;
    
    mac_send ether_send(
    .tx_go(tx_go),
    .rst_n(rst_n),
    .pyd_length(11'd46),   //payload�������ݳ���
        
    .src_mac(48'h00_0a_35_01_fe_c0),
    .des_mac(48'hFF_FF_FF_FF_FF_FF),
    .type_length(16'h08_06),
    
    .fifo_rdreq(fifo_rdreq),
    .fifo_rddata(fifo_rddata),
    .fifo_rdclk(fifo_rdclk),
        
    .crc_result(32'h69_1D_7D_96),
        
    .gmii_clk(gmii_clk),
    .gmii_tx_en(gmii_tx_en),
    .gmii_tx_err(gmii_tx_err),
    .gmii_tx_data(gmii_tx_data)
    );
            
    // ===========fifo���ݶ�ȡ==============
    reg [11:0] data_cnt;
    always@(posedge gmii_clk or negedge rst_n) begin
        if(!rst_n)
            data_cnt <= 12'd0;
        else if(fifo_rdreq)
            data_cnt <= data_cnt + 12'd1;
        else 
            data_cnt <= 12'd0;
    end
    
    // ��ȡarp�洢�����ֶΣ������ò��ұ���в���
    always@(*) begin
        case(data_cnt) 
            // ��̫��Э��
            0:fifo_rddata <= 8'h00;
            1:fifo_rddata <= 8'h01;
            
            // IPЭ��
            2:fifo_rddata <= 8'h08;
            3:fifo_rddata <= 8'h00;
            
            // MAC��ַ����
            4:fifo_rddata <= 8'h06;
            
            // IP��ַ����
            5:fifo_rddata <= 8'h04;
            
            // ������
            6:fifo_rddata <= 8'h00;
            7:fifo_rddata <= 8'h01;
            
            // ԴMAC��ַ
            8:fifo_rddata <= 8'h00;
            9:fifo_rddata <= 8'h0a;
            10:fifo_rddata <= 8'h35;
            11:fifo_rddata <= 8'h01;
            12:fifo_rddata <= 8'hfe;
            13:fifo_rddata <= 8'hc0;
            // ԴIP��ַ
            14:fifo_rddata <= 8'hC0;
            15:fifo_rddata <= 8'hA8;
            16:fifo_rddata <= 8'h00;
            17:fifo_rddata <= 8'h02;
            // Ŀ��MAC��ַ
            18:fifo_rddata <= 8'h00;
            19:fifo_rddata <= 8'h00;
            20:fifo_rddata <= 8'h00;
            21:fifo_rddata <= 8'h00;
            22:fifo_rddata <= 8'h00;
            23:fifo_rddata <= 8'h00;
            // Ŀ��IP��ַ
            24:fifo_rddata <= 8'hC0;
            25:fifo_rddata <= 8'hA8;
            26:fifo_rddata <= 8'h00;
            27:fifo_rddata <= 8'h03;
            // ����ֽ�
            28:fifo_rddata <= 8'h00;
            29:fifo_rddata <= 8'h00;
            30:fifo_rddata <= 8'hff;
            31:fifo_rddata <= 8'hff;
            32:fifo_rddata <= 8'hff;
            33:fifo_rddata <= 8'hff;
            34:fifo_rddata <= 8'hff;
            35:fifo_rddata <= 8'hff;
            36:fifo_rddata <= 8'h00;
            37:fifo_rddata <= 8'h23;
            38:fifo_rddata <= 8'hcd;
            39:fifo_rddata <= 8'h76;
            40:fifo_rddata <= 8'h63;
            41:fifo_rddata <= 8'h1a;
            42:fifo_rddata <= 8'h08;
            43:fifo_rddata <= 8'h06;
            44:fifo_rddata <= 8'h00;
            45:fifo_rddata <= 8'h01;
            default: fifo_rddata <= 8'h0;

        endcase
    
    end
         
    // ==========����֡���ͼ��================
    always@(posedge gmii_clk or negedge rst_n) begin
        if(!rst_n)
            cnt <= 25'd0;
        else
            cnt <= cnt + 25'd1;
    end
    
    assign tx_go = (cnt==1);
    
endmodule








