`timescale 1ns / 1ps

// ------------------------------------------------------------
// ��̫������ģ�飺�����л���ͬ��Э��
// ------------------------------------------------------------


module eth_ctrl(
    input                       clk,
    input                       rst,

    // ARP�˿��ź�
    input                       arp_rx_done         ,       // arp���Ľ������
    input                       arp_rx_type         ,       // arp���ձ������ͣ�0����1Ӧ��
    output     reg              arp_tx_en           ,       // arp����ʹ��
    output                      arp_tx_type         ,       // arp���ͱ������ͣ�0����1Ӧ��
    input                       arp_tx_done         ,       // arp���ͱ������
    input                       arp_gmii_tx_en      ,       // arp GMII���������Ч
    input               [7:0]   arp_gmii_txd        ,       // arp GMII��������

    // ICMP�˿��ź�
    input                       icmp_tx_start_en    ,       // icmp��ʼ�����ź�
    input                       icmp_tx_done        ,       // icmp��������ź�
    input                       icmp_gmii_tx_en     ,       // icmp GMII���������Ч�ź�
    input               [7:0]   icmp_gmii_txd       ,       // icmp GMII��������

    // GMII���ͽӿ�
    output                      gmii_tx_en          ,       // GMII���������Ч
    output              [7:0]   gmii_txd                    // GMII��������

    );

    // reg define
    reg         protocol_sw;                // Э���л��ź�
    reg         icmp_tx_busy;               // ICMP����æ״̬�ź�
    reg         arp_rx_flag;                // ���յ�ARP�����źű�־

    assign      arp_tx_type = 1'b1;         // �̶�arp��������ΪӦ��
    assign      gmii_tx_en  = protocol_sw ? icmp_gmii_tx_en : arp_gmii_tx_en;       // protocol_sw��0��arp���ģ�1��icmp����
    assign      gmii_txd    = protocol_sw ? icmp_gmii_txd : arp_gmii_txd;

    // ICMPæ�źſ���
    // always @(posedge clk or posedge rst) begin
    //     if(rst)
    //         icmp_tx_busy <= 1'b0;
    //     else if(icmp_tx_start_en)
    //         icmp_tx_busy <= 1'b1;
    //     else if(icmp_tx_done)
    //         icmp_tx_busy <= 1'b0;
    //     else;
    // end

    reg [23:0] icmp_timeout_cnt;  // 125MHzʱ��Լ0.134��

    always @(posedge clk or posedge rst) begin
        if (rst)
            icmp_timeout_cnt <= 0;
        else if (icmp_tx_start_en)
            icmp_timeout_cnt <= 0;
        else if (icmp_tx_busy && icmp_timeout_cnt < 24'hFFFFFF)
            icmp_timeout_cnt <= icmp_timeout_cnt + 1;
    end

    // �޸�icmp_tx_busy�߼�
    always @(posedge clk or posedge rst) begin
        if (rst)
            icmp_tx_busy <= 1'b0;
        else if (icmp_tx_start_en)
            icmp_tx_busy <= 1'b1;
        else if (icmp_tx_done || icmp_timeout_cnt == 24'hFFFFFF)  // ��ʱ��λ
            icmp_tx_busy <= 1'b0;
        else;
    end

    // ���ƽ��յ�ARP�����źű�־
    always @(posedge clk or posedge rst) begin
        if(rst)
            arp_rx_flag <= 1'b0;
        else if(arp_rx_done && (arp_rx_type == 1'b0))
            arp_rx_flag <= 1'b1;
        else
            arp_rx_flag <= 1'b0;
    end

    // ����protocol_sw�źź�arp_tx_en�ź�
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            protocol_sw <= 1'b0;
            arp_tx_en <= 1'b0;
        end
        else begin
            arp_tx_en <= 1'b0;
            if(icmp_tx_start_en) 
                protocol_sw <= 1'b1;
            else if(arp_rx_flag && (icmp_tx_busy == 1'b0)) begin
                protocol_sw <= 1'b0;
                arp_tx_en <= 1'b1;
            end
            else;
        end
    end

endmodule
