`timescale 1ns / 1ns

// -------------------------------------------------------
// arp testbench
// ͨ���Իػ�����arp�շ�
// -------------------------------------------------------

module tb_arp;

parameter T = 8;                                // ʱ������8ns
parameter OP_CYCLE = 100;                       // ��������

parameter  BOARD_MAC = 48'h00_11_22_33_44_55;        // �忨MAC��ַ
parameter  BOARD_IP  = {8'd192,8'd168,8'd0,8'd2}; 
// Ŀ��mac��ip
parameter  DES_MAC   = 48'hff_ff_ff_ff_ff_ff;
parameter  DES_IP  = {8'd192,8'd168,8'd0,8'd3}; 

// reg define
reg                 gmii_clk;
reg                 sys_rst;
reg                 arp_tx_en;
reg                 arp_tx_type;
reg     [3:0]       flow_cnt;
reg     [13:0]      delay_cnt;

// wire define
wire                gmii_rx_clk;
wire                gmii_rx_dv;
wire    [7:0]       gmii_rxd   ; //GMII��������
wire                gmii_tx_clk; //GMII����ʱ��
wire                gmii_tx_en ; //GMII��������ʹ���ź�
wire    [7:0]       gmii_txd   ; //GMII��������

wire                arp_rx_done; //ARP��������ź�
wire                arp_rx_type; //ARP�������� 0:����  1:Ӧ��
wire        [47:0]  src_mac    ; //���յ�Ŀ��MAC��ַ
wire        [31:0]  src_ip     ; //���յ�Ŀ��IP��ַ    
wire        [47:0]  des_mac    ; //���͵�Ŀ��MAC��ַ
wire        [31:0]  des_ip     ; //���͵�Ŀ��IP��ַ
wire                gmii_tx_done;
wire                arp_led;


assign  gmii_rx_clk = gmii_clk;
assign  gmii_tx_clk = gmii_clk;
assign  gmii_rx_dv  = gmii_tx_en;
assign  gmii_rxd    = gmii_txd;

assign  des_mac     = src_mac;
assign  des_ip      = src_ip;

initial begin
    gmii_clk        = 1'b0;
    sys_rst         = 1'b1;         // ��ʼ��λ
    #(T+1) sys_rst = 1'b0;
end

always #(T/2) gmii_clk = ~gmii_clk;

always @(posedge gmii_clk or posedge sys_rst) begin
    if(sys_rst) begin
        arp_tx_en <= 1'b0;
        arp_tx_type <= 1'b0;
        delay_cnt <= 1'b0;
        flow_cnt <= 1'b0;
    end
    else begin
        case (flow_cnt)
            4'd0 : flow_cnt <= flow_cnt + 4'd1;
            4'd1 : begin
                arp_tx_en <= 1'b1;
                arp_tx_type <= 1'b0;        // ����arp����
                flow_cnt <= flow_cnt + 4'd1;
            end
            4'd2 : begin
                arp_tx_en <= 1'b0;
                flow_cnt <= flow_cnt + 4'd1; 
            end
            4'd3 : begin
                if(gmii_tx_done) begin
                    flow_cnt <= flow_cnt + 4'd1;
                end
            end 
            4'd4 : begin
                delay_cnt <= delay_cnt + 14'd1;
                if(delay_cnt == OP_CYCLE - 1) begin
                    flow_cnt <= flow_cnt + 4'd1;
                end
            end
            4'd5 : begin
                arp_tx_en <= 1'b1;
                arp_tx_type <= 1'b1;        // arpӦ��
                flow_cnt <= flow_cnt + 4'd1;
            end
            4'd6 : begin
                arp_tx_en <= 1'b0;
                flow_cnt <= flow_cnt + 4'd1;
            end
            4'd7 : begin
                if(gmii_tx_done)
                    flow_cnt <= flow_cnt + 4'd1;
            end
            default:; 
        endcase
    end
end


// arpģ������
    arp #(
        .DES_IP             (DES_IP),
        .DES_MAC            (DES_MAC),
        .BOARD_IP           (BOARD_IP),
        .BOARD_MAC          (BOARD_MAC)
    )u_arp(
        .rst                (sys_rst),          
        .gmii_rx_clk        (gmii_rx_clk),
        .gmii_rx_dv         (gmii_rx_dv), 
        .gmii_rxd           (gmii_rxd),   
        .gmii_tx_clk        (gmii_tx_clk),
        .gmii_tx_en         (gmii_tx_en), 
        .gmii_txd           (gmii_txd),   
        .gmii_tx_done       (gmii_tx_done),          
        .arp_tx_en          (arp_tx_en),  
        .arp_tx_type        (arp_tx_type),
        .arp_rx_done        (arp_rx_done),
        .arp_rx_type        (arp_rx_type),
        .des_mac            (des_mac),    
        .des_ip             (des_ip),     
        .src_mac            (src_mac),    
        .src_ip             (src_ip),
        .arp_led            (arp_led)  
    );


endmodule
