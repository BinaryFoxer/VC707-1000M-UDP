`timescale 1ns / 1ps

// -------------------------------------------------------
// ��̫������Э�����ģ��
// ��ǰ֧��ARP��ICMP��UDP����Э���л�
// -------------------------------------------------------


module eth_ctrl_sw(
    input                   clk,
    input                   rst,

    // ARP�˿��ź�
    input                   arp_rx_done,                   // ARP���ݰ���������ź�
    input                   arp_rx_type,                   // ARP�������ͣ�0������1��Ӧ��
    output  reg             arp_tx_en,                     // ARP����ģ��ʹ���źţ���ʼ�����
    output                  arp_tx_type,                   // ARP�������ͣ�0������1��Ӧ��
    input                   arp_tx_done,                   // ARP�����������
    input                   arp_gmii_tx_en,                // ARPʹ��gmii_txd��������
    input           [7:0]   arp_gmii_txd,                  // ARPͨ��gmii_txd���͵�����

    // ICMP�˿��ź�
    input                   icmp_tx_start_en,              // ICMP����ģ��ʹ���źţ���ʼ�����
    input                   icmp_tx_done,                  // ICMP�����������
    input                   icmp_gmii_tx_en,               // ICMPʹ��gmii_txd��������
    input           [7:0]   icmp_gmii_txd,                 // ICMPͨ��gmii_txd���͵�����

    // ICMP fifo�ӿ��ź�
    input                   icmp_rec_en,                   // ICMP��������ʹ���ź�
    input           [7:0]   icmp_rec_data,
    input                   icmp_tx_req,                   // ICMP�����������ź�
    output          [7:0]   icmp_tx_data,                  // ICMP����������

    // UDP��ض˿��ź�
    input                   udp_tx_start_en,               // ICMP����ģ��ʹ���źţ���ʼ�����
    input                   udp_tx_done,                   // UDP��������ź�
    input                   udp_gmii_tx_en,                // UDPʹ��gmii_txd��������
    input           [7:0]   udp_gmii_txd,                  // UDPͨ��gmii_txd���͵�����

    // UDP fifo�ӿ��ź�
    input                   udp_rec_en,                   // ICMP��������ʹ���ź�
    input           [7:0]   udp_rec_data,
    input                   udp_tx_req,                   // ICMP�����������ź�
    output          [7:0]   udp_tx_data,                  // ICMP����������

    // fifo�ӿ��ź�
    input           [7:0]   tx_data,                      // ����������
    output                  tx_req,
    output  reg             rec_en,
    output  reg     [7:0]   rec_data,

    // GMII��������
    output  reg             gmii_tx_en,
    output  reg     [7:0]   gmii_txd
    );

    // define reg
    reg [1:0]   protocol_sw;
    reg         icmp_tx_busy;
    reg         udp_tx_busy;
    reg         arp_rx_flag;
    reg         icmp_tx_req_d0;
    reg         udp_tx_req_d0;

    assign  arp_tx_type = 1'b1;                         // �����ã�ֻ��Ӧ��
    assign  tx_req = udp_tx_req ? 1'b1 : icmp_tx_req;
    assign  icmp_tx_data = icmp_tx_req_d0 ? tx_data : 8'd0;
    assign  udp_tx_data = udp_tx_req_d0 ? tx_data : 8'd0;

    // �Ĵ�һ�������źţ�������������һ��
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            icmp_tx_req_d0 <= 1'b0;
            udp_tx_req_d0 <= 1'b0;
        end
        else begin
            icmp_tx_req_d0 <= icmp_tx_req;
            udp_tx_req_d0 <= udp_tx_req;
        end
    end

    // ����ʹ���ź��жϽ�������
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            rec_en  <= 1'b0;
            rec_data <= 8'd0;
        end
        else if(icmp_rec_en) begin
            rec_en <= icmp_rec_en;
            rec_data <= icmp_rec_data;
        end
        else if(udp_rec_en) begin
            rec_en <= udp_rec_en;
            rec_data <= udp_rec_data;
        end
        else begin
            rec_en <= 1'b0;
            rec_data <= rec_data;
        end
    end

    // Э���л�
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            gmii_tx_en <= 1'b0;
            gmii_txd <= 8'd0;
        end
        else begin
            case(protocol_sw)
                2'b00:begin
                    gmii_tx_en <= arp_gmii_tx_en;
                    gmii_txd   <= arp_gmii_txd;
                end

                2'b01:begin
                    gmii_tx_en <= icmp_gmii_tx_en;
                    gmii_txd   <= icmp_gmii_txd;
                end

                2'b10:begin
                    gmii_tx_en <= udp_gmii_tx_en;
                    gmii_txd   <= udp_gmii_txd;
                end

                default: ;
            endcase
        end
    end

    // ��ʱ�������
    reg [23:0] timeout_cnt;  // 125MHzʱ��Լ0.134��

    always @(posedge clk or posedge rst) begin
        if (rst)
            timeout_cnt <= 0;
        else if (icmp_tx_start_en)
            timeout_cnt <= 0;
        else if ((icmp_tx_busy && timeout_cnt < 24'hFFFFFF) || (udp_tx_busy && timeout_cnt < 24'hFFFFFF))
            timeout_cnt <= timeout_cnt + 1;
    end


    // ����ICMP����æ�ź�
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            icmp_tx_busy <= 1'b0;
        end
        else if(icmp_tx_start_en) begin
            icmp_tx_busy <= 1'b1;
        end
        else if(icmp_tx_done || timeout_cnt == 24'hFFFFFF) begin
            icmp_tx_busy <= 1'b0;
        end
        else;
    end

    // ����UDP����æ�ź�
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            udp_tx_busy <= 1'b0;
        end
        else if(udp_tx_start_en) begin
            udp_tx_busy <= 1'b1;
        end
        else if(udp_tx_done || timeout_cnt == 24'hFFFFFF) begin
            udp_tx_busy <= 1'b0;
        end
        else;
    end

    // ����ARP���������־
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            arp_rx_flag <= 1'b0;
        end
        else if(arp_rx_done && (arp_rx_type == 1'b0))
            arp_rx_flag <= 1'b1;
        else 
            arp_rx_flag <= 1'b0;
    end

    // ����protocolЭ���л��źź�arp_tx_en�ź�
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            protocol_sw <= 2'b00;
            arp_tx_en   <= 1'b0;
        end
        else begin
            arp_tx_en <= 1'b0;
            if(udp_tx_start_en)
                protocol_sw <= 2'b10;
            else if(icmp_gmii_tx_en)
                protocol_sw <= 2'b01;
            else if((arp_rx_flag && (udp_tx_busy == 1'b0)) || (arp_rx_flag && (icmp_tx_busy == 1'b0))) begin
                protocol_sw <= 2'b00;
                arp_tx_en <= 1'b1;
            end
            else;
        end
    end


endmodule
