`timescale 1ns / 1ps

// -----------------------------------
// arp����ģ��
// -----------------------------------

module arp(
    input               rst,
    // gmii�ӿ�
    input               gmii_rx_clk,                    // gmii����ʱ��
    input               gmii_rx_dv,                     // gmii����������Ч
    input        [7:0]  gmii_rxd,                       // gmii��������
    input               gmii_tx_clk,                    // gmii����ʱ��
    output              gmii_tx_en,                     // gmii����ʹ��
    output       [7:0]  gmii_txd,                       // gmii��������
    output              gmii_tx_done,                   // ��̫���������

    // �û��ӿ�
    input               arp_tx_en,                      // arp����ʹ��
    input               arp_tx_type,                    // ����arp��֡���ͣ�0����1Ӧ��
    output              arp_rx_done,                    // arp�����������
    output              arp_rx_type,                    // ����arp֡���ͣ�0����1Ӧ��
    input        [47:0] des_mac,                        // Ŀ��mac��ַ
    input        [31:0] des_ip,                         // Ŀ��ip
    output       [47:0] src_mac,                        // Դmac��ַ
    output       [31:0] src_ip                           // Դip��ַ
    );

    // parameter define
    // �忨mac��ip
    parameter BOARD_MAC = 48'h00_0a_35_01_fe_c0;        // �忨MAC��ַ
    parameter BOARD_IP  = 32'hC0_A8_00_02;              // �忨IP��ַ
    // Ŀ��mac��ip
    parameter   DES_MAC   = 48'hA8_2B_DD_25_DA_43;      // PC mac
    parameter   DES_IP    = 32'hC0_A8_00_03;            // PC ip

    // wire define
    wire          crc_en;             // crc��ʼ��������ʹ��
    wire          crc_clr;            // crc��λ�ź�
    wire   [7:0]  data;               // ����У���8λ����
    wire  [31:0]  crc_data;           // CRCУ������
    wire  [31:0]  crc_next;           // �´�У�������CRC����

    assign  data = gmii_txd;

    arp_tx #(
        .BOARD_IP(BOARD_IP),
        .BOARD_MAC(BOARD_MAC),
        .DES_IP(DES_IP),
        .DES_MAC(DES_MAC)
    ) u_arp_tx(
        .clk(gmii_tx_clk),        
        .rst(rst),        
        .arp_tx_en(arp_tx_en),  
        .arp_tx_type(arp_tx_type),
        .des_mac(des_mac),    
        .des_ip(des_ip),     
        .crc_data(crc_data),   
        .crc_next(crc_next[31:24]),   
        .crc_en(crc_en),     
        .crc_clr(crc_clr),    
        .gmii_txd(gmii_txd),   
        .gmii_tx_en(gmii_tx_en), 
        .gmii_tx_done(gmii_tx_done)
    );

    arp_rx #(
        .BOARD_IP(BOARD_IP),
        .BOARD_MAC(BOARD_MAC)
    )u_arp_rx(
        .rst(rst),       
        .clk(gmii_rx_clk),                   
        .gmii_rx_dv(gmii_rx_dv),
        .gmii_rxd(gmii_rxd),           
        .arp_rx_done(arp_rx_done),
        .arp_rx_type(arp_rx_type),
        .src_ip(src_ip),    
        .src_mac(src_mac)    

    );

    CRC32_d8 u_crc32_d8(
        .clk(gmii_tx_clk),    
        .rst(rst),    
        .crc_en(crc_en), 
        .crc_clr(crc_clr),
        .data(data),        
        .crc_data(crc_data),
        .crc_next(crc_next)
    );

endmodule
