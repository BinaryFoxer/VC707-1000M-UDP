`timescale 1ns / 1ps

// -----------------------------------------------------------------
// arp����ģ��,ͨ��arpģ�鷢������
// -----------------------------------------------------------------


module arp_ctrl(
    input               clk,
    input               sys_rst,

    input               touch_key,                  // ����������������arp����
    input               arp_rx_done,                // ARP�����������
    input               arp_rx_type,                // ARP�������� 0:����  1:Ӧ�� 
    output   reg        arp_tx_en,                  // ARP����ʹ��
    output   reg        arp_tx_type                 // ARP�������� 0:����  1:Ӧ��
    );

    // reg define
    reg             touch_key_d0;
    reg             touch_key_d1;

    // wire define
    wire            pos_touch_key;

    assign pos_touch_key = ~touch_key_d1 & touch_key_d0;

    // ��ʱ������touch_key�źŲɼ�������
    always @(posedge clk or posedge sys_rst) begin
        if(sys_rst) begin
            touch_key_d0 <= 1'b0;
            touch_key_d1 <= 1'b0;
        end
        else begin
            touch_key_d0 <= touch_key;
            touch_key_d1 <= touch_key_d0;
        end
    end

    // ��ֵ��arp���ͺ�arp����
    always @(posedge clk or posedge sys_rst) begin
        if(sys_rst) begin
            arp_tx_en <= 1'b0;
            arp_tx_type <= 1'b0;
        end
        else begin
            if(pos_touch_key) begin
                arp_tx_en <= 1'b1;                  // ����arpʹ��
                arp_tx_type <= 1'b0;                // ����arp����
            end
            else if((arp_rx_done == 1'b1) && (arp_tx_type == 1'b0)) begin   // ���յ�arp����,����arpӦ��
                arp_tx_en <= 1'b1;
                arp_tx_type <= 1'b1;
            end
            else 
                arp_tx_en <= 1'b0;
        end
    end

endmodule
